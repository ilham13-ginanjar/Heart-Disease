��      �sklearn.ensemble._forest��RandomForestClassifier���)��}�(�base_estimator��sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �_sklearn_version��1.0.2�ub�n_estimators�Kd�estimator_params�(hhhhhhhhhht��	bootstrap���	oob_score���n_jobs�J����hK*�verbose�K �
warm_start��hN�max_samples�NhhhKhKhKhG        h�auto�hNhG        hG        �feature_names_in_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h)�dtype����O8�����R�(K�|�NNNJ����J����K?t�b�]�(�age��sex��cp��trestbps��chol��fbs��restecg��thalach��exang��oldpeak��slope��ca��thal�et�b�n_features_in_�K�
n_outputs_�K�classes_�h(h+K ��h-��R�(KK��h2�i8�����R�(K�<�NNNJ����J����K t�b�C               �t�b�
n_classes_�K�base_estimator_�h	�estimators_�]�(h)��}�(hhhhhKhKhKhG        hh$hNhJf��_hG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��h2�f8�����R�(KhQNNNJ����J����K t�b�C              �?�t�bhUh&�scalar���hPC       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���Kh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hK�
node_count�K1�nodes�h(h+K ��h-��R�(KK1��h2�V56�����R�(Kh6N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(h�h2�i8�����R�(KhQNNNJ����J����K t�bK ��h�h�K��h�h�K��h�haK��h�haK ��h�h�K(��h�haK0��uK8KKt�b�B�
                             �?�>$�*��?�           8�@                           @B�b-jX�?�            �w@                           �?`RC4%�?�             q@                          �T@T�����?�            �l@������������������������       �                     �?                          �c@l�b�G��?�            �l@������������������������       �      �?�             l@������������������������       �      �?             @	                          �b@v ��?            �E@
                          �h@������?             ;@������������������������       �                     &@������������������������       �     ��?
             0@������������������������       �                     0@                          �c@�q�q�?F            �[@                          8p@� ���?3            @S@                           �?d}h���?             E@������������������������       �������?            �B@������������������������       �                     @                           �?�#-���?            �A@������������������������       ��z�G��?             $@������������������������       �                     9@                           l@�������?             A@������������������������       �                     *@                           �?և���X�?             5@������������������������       ��<ݚ�?             "@������������������������       �r�q��?             (@       $                    �?�^��T��?�             m@       #                    @^n����?)             N@                           �s@ZՏ�m|�?             �H@              	          033@�Ra����?             F@������������������������       ��(\����?             D@������������������������       �                     @!       "                    w@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �        	             &@%       *                    �?&^�)b�?w            �e@&       )                    `@@;�"�?Q            �^@'       (                    �L@t�U����?+            �P@������������������������       �                    �@@������������������������       �������?             A@������������������������       �        &             L@+       .       
             �?�`���?&            �H@,       -       	          ����?�LQ�1	�?             7@������������������������       �      �?             @������������������������       �                     3@/       0       	          hff@���B���?             :@������������������������       �      �?             8@������������������������       �                      @�t�b�values�h(h+K ��h-��R�(KK1KK��ha�B       �p@     �u@     �[@      q@     �B@     `m@      1@     �j@      �?              0@     �j@      ,@     @j@       @       @      4@      7@      4@      @      &@              "@      @              0@     �R@     �B@     @P@      (@     �@@      "@     �@@      @              @      @@      @      @      @      9@              "@      9@              *@      "@      (@      @       @       @      $@     �c@     @R@      3@     �D@       @     �D@      @     �C@      �?     �C@      @              @       @      @                       @      &@             �a@      @@     �\@       @     �M@       @     �@@              :@       @      L@              9@      8@      4@      @      �?      @      3@              @      5@      @      5@       @        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ�=�KhG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK/hyh(h+K ��h-��R�(KK/��h��BH
                             �?;�׊��?�           8�@                           �?�š�9�?�            �v@                           q@�'F����?�            �o@                           �N@8EGr��?}             i@                           �M@ �<#�?n            �e@������������������������       �������?g            �d@������������������������       ��eP*L��?             &@������������������������       �                     9@	              	          033�?�q�q�?!             K@
              	          ����? �o_��?             I@������������������������       �     ��?             @@������������������������       �        
             2@������������������������       �                     @                           @^H���+�?B            �[@                           �?�q�q�?             H@              	          `ff�?X�Cc�?             ,@������������������������       �                     @������������������������       �                     "@                           �?��hJ,�?             A@������������������������       �     ��?	             0@������������������������       �                     2@              
             �?�[|x��?&            �O@                           �?���J��?            �I@������������������������       �                    �F@������������������������       �r�q��?             @                           `@�q�q�?             (@������������������������       �                     @������������������������       �և���X�?             @       &                    �?������?�            @o@                           �E@�F}ʽx�?`            �b@������������������������       �        	             *@        #                    �?�q�q�?W            @a@!       "                    �?r�qG�?             H@������������������������       �`�Q��?             9@������������������������       �                     7@$       %                    @r�q��?:            �V@������������������������       ����tT��?7            �U@������������������������       �                     @'       (                   @X@���F6��?D            �X@������������������������       �                     �?)       ,       	          ����?��<D�m�?C            �X@*       +       	          833�?PN��T'�?             ;@������������������������       � �q�q�?             8@������������������������       �                     @-       .       
             �?�J�T�?3            �Q@������������������������       �        /            �P@������������������������       ����Q��?             @�t�bh�h(h+K ��h-��R�(KK/KK��ha�B�       �r@     �s@      \@     �o@      D@     �j@      6@     @f@      6@      c@      0@     �b@      @      @              9@      2@      B@      ,@      B@      ,@      2@              2@      @              R@     �C@      ,@      A@      "@      @              @      "@              @      =@      @      &@              2@      M@      @      I@      �?     �F@              @      �?       @      @      @              @      @      g@     �P@      W@     �M@              *@      W@      G@      1@      ?@      1@       @              7@     �R@      .@     �R@      &@              @      W@      @              �?      W@      @      7@      @      7@      �?              @     @Q@       @     �P@              @       @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ\bshG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK1hyh(h+K ��h-��R�(KK1��h��B�
                            Pb@�p ��?~           8�@                           �?��h��?�            �p@                          @\@�Q����?H             ^@                            G@؇���X�?             <@                          �`@���Q��?             $@������������������������       ��q�q�?             @������������������������       �                     @������������������������       �                     2@	                          m@n>�X�q�?7             W@
                          �]@��S���?            �F@������������������������       �                      @������������������������       ���J�fj�?            �B@              
             �?�*/�8V�?            �G@������������������������       �z�G�z�?             @������������������������       ���s����?             E@              	          ����?��"Ҥ(�?b            �b@                          �p@�2�IQ�?9            �V@                           @����0�?"             K@������������������������       �����X�?            �H@������������������������       �                     @������������������������       �                     B@������������������������       �        )            �N@       $                    �?���$�?�            �u@              	          033@�3d`��?�            �k@                           @��UV�?�            �j@                           @N@p��D׀�?`            �c@������������������������       � �}�$>�?U            �a@������������������������       ���S���?             .@                           �?��N`.�?!            �K@������������������������       ��5��?             ;@������������������������       �@4և���?             <@        #                    @և���X�?             @!       "                    @J@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @%       *                   �k@�U���?M             _@&       '                   �d@�GN�z�?             6@������������������������       �                      @(       )                   p`@R���Q�?             4@������������������������       �      �?             @������������������������       �        
             ,@+       .                    �?�!���?=            �Y@,       -                    @�GN�z�?(            �P@������������������������       �և���X�?            �A@������������������������       �                     ?@/       0                   `c@      �?             B@������������������������       �                     $@������������������������       ��	j*D�?             :@�t�bh�h(h+K ��h-��R�(KK1KK��ha�B       �r@     �s@     `h@      S@     �O@     �L@      @      8@      @      @      @       @              @              2@     �M@     �@@      8@      5@       @              0@      5@     �A@      (@      �?      @      A@       @     �`@      3@     �Q@      3@     �A@      3@     �A@      ,@              @      B@             �N@             @Z@     �m@      ?@     �g@      ;@     @g@      "@     �b@       @     �a@      @       @      2@     �B@      0@      &@       @      :@      @      @       @      @              @       @               @             �R@      I@      @      1@       @              @      1@      @      @              ,@     @Q@     �@@     �I@      .@      4@      .@      ?@              2@      2@              $@      2@       @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ��.hG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK3hyh(h+K ��h-��R�(KK3��h��B(                            pb@��FY��?�           8�@                           @�lr�]��?�            �p@                           �?l��[B��?L             ]@                          pr@4և����?&             L@                           �G@r�����?#            �J@������������������������       ����Q��?	             .@������������������������       ��KM�]�?             C@������������������������       �                     @	              
             �?d��0u��?&             N@
                          �r@ �q�q�?             H@������������������������       � qP��B�?            �E@������������������������       �z�G�z�?             @                          �j@�8��8��?             (@������������������������       �                     �?������������������������       �                     &@              	          833�?f�8A_�?]            �b@                          �a@�5��?             ;@                           �L@8����?             7@������������������������       ����|���?	             &@������������������������       �                     (@������������������������       �                     @                           �?`Jj��?K             _@������������������������       �        A             [@                           �O@      �?
             0@������������������������       ����!pc�?             &@������������������������       �                     @       (                    �?����S��?�            �u@       #                    @L�A���?[             b@                            �?�~�4_��?9             V@                           �L@��ɉ�?)            @P@������������������������       �                     F@������������������������       �և���X�?             5@!       "       	             �?\X��t�?             7@������������������������       �j���� �?             1@������������������������       �                     @$       '                   �n@l�b�G��?"            �L@%       &       
             �?\-��p�?             =@������������������������       �                     "@������������������������       �z�G�z�?             4@������������������������       �                     <@)       .                    �?��9~��?|            `i@*       +                    @G@x̓��s�?l            �e@������������������������       �        -            �R@,       -                    @Ș����??             Y@������������������������       ���(\���?3             T@������������������������       ��G�z��?             4@/       2                    �?���>4��?             <@0       1                    _@     ��?	             0@������������������������       �և���X�?             @������������������������       �                     "@������������������������       �                     (@�t�bh�h(h+K ��h-��R�(KK3KK��ha�B0       r@     `t@     `g@      T@      N@      L@      *@     �E@      $@     �E@      @      "@      @      A@      @             �G@      *@      G@       @      E@      �?      @      �?      �?      &@      �?                      &@     �_@      8@      &@      0@      @      0@      @      @              (@      @              ]@       @      [@               @       @      @       @      @             �Y@     �n@      R@     @R@      3@     @Q@      "@      L@              F@      "@      (@      $@      *@      $@      @              @     �J@      @      9@      @      "@              0@      @      <@              >@     �e@      1@     �c@             �R@      1@     �T@      @     �R@      &@      "@      *@      .@      *@      @      @      @      "@                      (@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJj�c;hG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK7hyh(h+K ��h-��R�(KK7��h��B                             @|��z��?�           8�@                           �?6�Զ�?�             w@       
       
             �?�Uo���?]             c@                           �?8^s]e�?5            �U@              	          033�?�n_Y�K�?            �C@������������������������       ���a�n`�?             ?@������������������������       �                      @       	                    �?      �?             H@������������������������       �z�G�z�?	             .@������������������������       �                    �@@                            P@�θ�?(            @P@                          xt@�t����?             �I@������������������������       �t��ճC�?             F@������������������������       �և���X�?             @                           �?X�Cc�?             ,@������������������������       �      �?              @������������������������       �                     @                           �?�~i��?�            @k@                          �m@�r�MȢ?A            �Z@                           �K@`'�J�?            �I@������������������������       �                    �D@������������������������       �z�G�z�?             $@������������������������       �        $             L@                           c@���GYW�?M            �[@              	          ����?l��w��?G            �Y@������������������������       �0�,���?-            �P@������������������������       �b�2�tk�?             B@                           m@      �?              @������������������������       �                     @������������������������       �      �?             @       *       
             �?4�2%ޑ�?�            �n@        %                   �d@fP*L���?k             f@!       $                   �g@�����H�?\             c@"       #                    @tX�}}��?Z            �b@������������������������       � 	��p�?W             b@������������������������       �r�q��?             @������������������������       �                      @&       '                    @\X��t�?             7@������������������������       �                     (@(       )       
             �?�C��2(�?             &@������������������������       �                     @������������������������       �؇���X�?             @+       2                   �^@���=�/�?-            @Q@,       /                    �?�GN�z�?             6@-       .       	          833�?      �?	             0@������������������������       ���S�ۿ?             .@������������������������       �                     �?0       1       	          ����?      �?             @������������������������       �                      @������������������������       �      �?             @3       4                    i@�*/�8V�?             �G@������������������������       �                     @5       6                    �?r�q��?             E@������������������������       �l��\��?             A@������������������������       �      �?              @�t�bh�h(h+K ��h-��R�(KK7KK��ha�Bp        r@     pt@     �X@     �p@     �R@     @S@      N@      ;@      .@      8@      @      8@       @             �F@      @      (@      @     �@@              .@      I@      @     �F@      @     �D@      @      @      "@      @      @      @      @              8@     @h@       @     @Z@       @     �H@             �D@       @       @              L@      6@     @V@      0@     �U@       @     @P@      ,@      6@      @       @      @               @       @     �g@      L@     �b@      ;@      a@      1@      a@      .@     �`@      $@      �?      @               @      *@      $@      (@              �?      $@              @      �?      @      D@      =@      @      1@       @      ,@      �?      ,@      �?              @      @               @      @      �?     �A@      (@              @     �A@      @      ?@      @      @      @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJGԙGhG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK#hyh(h+K ��h-��R�(KK#��h��B�                             �?�������?�           8�@                          0f@�	4!���?�            pq@       
                    �Q@�����?�            �p@                           �?J���?�            pp@              
             �?և���X�?=            �V@������������������������       ��GN�z�?              F@������������������������       �֭��F?�?            �G@       	                    �?Du9iH��?m            �e@������������������������       ��䞠�l�?0            @S@������������������������       ��==Q�P�?=            �W@                           �?�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     $@                           @�\`*��?�             u@                           @�K<��V�?�            �r@                           �?��M[�?�             k@              
             �?�YX�Z�?d            �d@������������������������       ��r����?            �F@������������������������       ���v$���?H            �^@                           �?~���L0�?%            �H@������������������������       �                     @������������������������       ���s����?             E@              	          `ff�?�p ��?0            �T@                          �a@�Z4���?)            �P@������������������������       ��<ݚ�?	             2@������������������������       ����c�H�?             �H@������������������������       �                     .@                          �l@D�n�3�?             C@������������������������       �        	             *@               
             �?��H�}�?             9@������������������������       �                     @!       "                    �?���N8�?             5@������������������������       �@4և���?             ,@������������������������       �և���X�?             @�t�bh�h(h+K ��h-��R�(KK#KK��ha�B0       Pr@      t@     �j@     @P@     �j@     �K@     �j@     �I@      J@     �C@      A@      $@      2@      =@      d@      (@      Q@      "@      W@      @       @      @              @       @                      $@     �S@     p@     �O@     `m@      7@      h@       @     �c@      @     �C@       @      ^@      .@      A@      @               @      A@      D@      E@      9@      E@      ,@      @      &@      C@      .@              0@      6@              *@      0@      "@              @      0@      @      *@      �?      @      @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ��AhG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK/hyh(h+K ��h-��R�(KK/��h��BH
                            �b@�������?�           8�@       	                   �\@�)!�,�?�            �r@                          pj@0,Tg��?             E@������������������������       �                     5@                           �?�G��l��?             5@������������������������       �                     "@                          �l@�8��8��?             (@������������������������       �z�G�z�?             @������������������������       �                     @
                           �?�R��Hx�?�             p@                           �F@�d����?E            �^@                            D@�����H�?             "@������������������������       �                     �?������������������������       �                      @                          0`@�q�q�??            �\@������������������������       �t/*�?            �G@������������������������       ���:c���?'            �P@              	          ����?��S�ۿ?Q            �`@                          @]@ҳ�wY;�?             1@������������������������       �                     @������������������������       �                     &@                          pb@���<_�?F            �]@������������������������       ��L��ȕ?7            @W@������������������������       �HP�s��?             9@       $                    @��c���?�            �s@                           @L@�L����?�            @o@                           �?H�!b	�?j            @d@              	          ����?BӀN��?b            �b@������������������������       �|)����?;            �V@������������������������       �        '             N@������������������������       �                     &@        #       	          033@      �?4             V@!       "                    a@<�\`*��?0             U@������������������������       �և���X�?            �A@������������������������       �Jm_!'1�?            �H@������������������������       �                     @%       *                    �?�G\�c�?3            @P@&       )                    �?>A�F<�?             C@'       (                    @K@b�2�tk�?             2@������������������������       �������?             .@������������������������       �                     @������������������������       �                     4@+       .                   �q@������?             ;@,       -       	          hff @r�q��?             8@������������������������       �                     4@������������������������       �                     @������������������������       �                     @�t�bh�h(h+K ��h-��R�(KK/KK��ha�B�       Pr@      t@     �j@     �U@      &@      ?@              5@      &@      $@              "@      &@      �?      @      �?      @             `i@     �K@     @S@      G@      �?       @      �?                       @      S@      C@     �C@       @     �B@      >@     �_@      "@      &@      @              @      &@             �\@      @      W@      �?      7@       @     �S@     �m@     �D@      j@       @     @c@       @     �a@       @     �T@              N@              &@     �@@     �K@      =@     �K@      4@      .@      "@      D@      @              C@      ;@      ?@      @      &@      @      &@      @              @      4@              @      4@      @      4@              4@      @              @        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ,�hG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK-hyh(h+K ��h-��R�(KK-��h��B�	                             �?&n.���?�           8�@       	                   `b@М��O�?}            �g@                           �?����*��?(            �M@                          �`@�	j*D�?            �C@                           @�q�q�?             2@������������������������       �$�q-�?
             *@������������������������       �                     @������������������������       �                     5@������������������������       �                     4@
                           @L@��2(&�?U            �`@������������������������       �        1             S@              	          `ff�?��X��?$             L@                           �N@:	��ʵ�?            �F@������������������������       �և���X�?             ,@������������������������       �                     ?@                          c@�C��2(�?             &@������������������������       �                     �?������������������������       �                     $@                            �?�J����?	           �z@              	          pff�?��V#�?�            �j@                           �?�F�j��?@            �Z@                          �e@��f/w�?$            �N@������������������������       ��G�z�?             D@������������������������       �                     5@                           �?�r����?            �F@������������������������       �@�0�!��?             A@������������������������       �                     &@              	           33@>����?D            @[@                            J@(N:!���?A            @Z@������������������������       �      �?             8@������������������������       � 7���B�?3            @T@������������������������       �                     @!       (       	          ����?�g\Ɋ�?�             j@"       %                    �?p�}�ޤ�?b            @b@#       $                    @     ��?B             X@������������������������       �`���i��?>             V@������������������������       �      �?              @&       '                    �?���H.�?              I@������������������������       �4���C�?            �@@������������������������       ��t����?             1@)       *                    �B@؇���X�?#            �O@������������������������       �                      @+       ,                    �?Xny��?"            �N@������������������������       � �o_��?             9@������������������������       �                     B@�t�bh�h(h+K ��h-��R�(KK-KK��ha�B�       �q@     �t@     �F@     @b@      ;@      @@      ;@      (@      @      (@      �?      (@      @              5@                      4@      2@     �\@              S@      2@      C@       @     �B@       @      @              ?@      $@      �?              �?      $@             �m@     `g@      b@     �Q@      J@      K@      *@      H@      *@      ;@              5@     �C@      @      <@      @      &@             @W@      0@     @W@      (@      .@      "@     �S@      @              @      W@     @]@      C@      [@      "@     �U@      @     @T@       @      @      =@      5@      ,@      3@      .@       @      K@      "@               @      K@      @      2@      @      B@        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJf��'hG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK/hyh(h+K ��h-��R�(KK/��h��BH
                             �?JGC8{��?�           8�@                           @2\Q��?           Py@       
                    �?�����?�            pq@                           �?`.��A��?�            �m@                          �s@����q�?I            @[@������������������������       �        A            @X@������������������������       �r�q��?             (@       	                    �?��ɉ�?R            @`@������������������������       �z�G�z�?#            �K@������������������������       ����Lͩ�?/            �R@                          hs@�Q����?             D@                           d@�ʻ����?             A@������������������������       ��q�q�?             5@������������������������       �$�q-�?             *@������������������������       �                     @              	          ����?����1�?R            �_@                          �c@����e��?,            �P@                          c@�<ݚ�?             B@������������������������       ��q�q�?             5@������������������������       ���S�ۿ?             .@                           �?���Q��?             >@������������������������       �����X�?             ,@������������������������       �      �?
             0@                          pe@d��0u��?&             N@              
             �?�:�]��?#            �I@������������������������       ��Ń��̧?             E@������������������������       ��q�q�?             "@������������������������       �                     "@       $                   �b@�϶O'3�?�            @j@       #                   �p@dOwq=)�?n             e@                           �Z@Ș����?D             Y@������������������������       �                     @!       "                    @N@�j�@�?@            �W@������������������������       ���ɉ�?-            @P@������������������������       ��q�q�?             >@������������������������       �        *            @Q@%       *                    �M@#z�i��?            �D@&       '                    �D@������?             A@������������������������       �                     @(       )       	          ���@�r����?             >@������������������������       �@4և���?             <@������������������������       �                      @+       ,                    �O@؇���X�?             @������������������������       �                     @-       .                    �?�q�q�?             @������������������������       �                     �?������������������������       �      �?              @�t�bh�h(h+K ��h-��R�(KK/KK��ha�B�       �q@     �t@     �\@     0r@     �D@     �m@      4@     `k@       @     �Z@             @X@       @      $@      2@      \@      &@      F@      @      Q@      5@      3@      .@      3@      ,@      @      �?      (@      @             @R@     �J@      :@      D@       @      <@      @      ,@      �?      ,@      2@      (@      @      $@      ,@       @     �G@      *@     �G@      @     �D@      �?      @      @              "@     �d@      F@      c@      1@     �T@      1@              @     �T@      (@     �O@       @      4@      $@     @Q@              ,@      ;@       @      :@      @              @      :@       @      :@       @              @      �?      @               @      �?      �?              �?      �?�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJy"rhG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK7hyh(h+K ��h-��R�(KK7��h��B                	             �?Z�����?�           8�@                           �?*t�*�N�?�            �r@       
                    �?JJ����?D            �W@                           @t�F�}�?%            �I@                          xt@r�q��?             B@������������������������       �<���D�?            �@@������������������������       ��q�q�?             @       	                   �c@��S���?             .@������������������������       �r�q��?             @������������������������       ��q�q�?             "@                          @[@�^�����?            �E@                           �?      �?              @������������������������       �                     �?������������������������       �                     @              	          833�?b�h�d.�?            �A@������������������������       � 	��p�?             =@������������������������       ��q�q�?             @                           �K@�d2 Λ�?�            �i@                           @hA� �?W            �a@                          @[@@���a��?J            �\@������������������������       �      �?              @������������������������       �        C            �Z@                          Pd@z�G�z�?             9@������������������������       �        
             3@������������������������       �r�q��?             @                          �l@     ��?)             P@������������������������       �                     8@                           �?H�z�G�?             D@������������������������       �ҳ�wY;�?
             1@������������������������       ���+7��?             7@       *                   pb@J�WrV�?�            �s@        %                    �?*K�U��?�            `j@!       "                    i@j���� �?             A@������������������������       �                     @#       $                    �?����X�?             <@������������������������       ����N8�?             5@������������������������       �                     @&       '                    @I@N�hƇ�?j             f@������������������������       �                    �F@(       )                    �?�禺f��?P            �`@������������������������       �*;L]n�?             >@������������������������       ����J��?=            �Y@+       2                   �l@�ǧ\�?F            �Z@,       /                    �?h�����?#             L@-       .       	          033�?�q�q�?             B@������������������������       �                     @������������������������       ���a�n`�?             ?@0       1                   Pi@P���Q�?             4@������������������������       �                     �?������������������������       �                     3@3       4                    @z�G�z�?#             I@������������������������       �                     >@5       6                   �_@      �?             4@������������������������       �                     @������������������������       �����X�?             ,@�t�bh�h(h+K ��h-��R�(KK7KK��ha�Bp       �q@     �t@     �P@     �l@      F@      I@      ,@     �B@      @      >@      @      =@       @      �?       @      @      @      �?      @      @      >@      *@      �?      @      �?                      @      =@      @      ;@       @       @      @      7@     �f@      @     �`@      �?     �\@      �?      @             �Z@      @      4@              3@      @      �?      1@     �G@              8@      1@      7@      &@      @      @      1@     `k@     �X@     @f@     �@@      4@      ,@              @      4@       @      4@      �?              @     �c@      3@     �F@             @\@      3@      *@      1@      Y@       @     �D@     @P@      ?@      9@      (@      8@      @              @      8@      3@      �?              �?      3@              $@      D@              >@      $@      $@              @      $@      @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ�A�'hG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK1hyh(h+K ��h-��R�(KK1��h��B�
                             @K@V���Ş�?�           8�@                           @� Ђ���?�            �r@                           �?���L���?�            @k@              	          `ff@`Jj��?q            @g@                          �]@�.ߴ#�?p            �f@������������������������       �r�q��?"             K@������������������������       �        N             `@������������������������       �                     @	              	          ����?     ��?             @@
                           ]@�㙢�c�?             7@������������������������       �                     @������������������������       �                     3@������������������������       �                     "@                          0b@��i#[�?6             U@������������������������       �                     @@                          �^@      �?!             J@                           �D@z�G�z�?             9@������������������������       �                     @������������������������       ��C��2(�?             6@              	             �?�<ݚ�?             ;@������������������������       �        
             2@������������������������       ��q�q�?             "@       &       	          ����?*܂��q�?�            �s@                           l@༉p���?�            �j@                           �?     ��?(             P@              	          pff�?8��8���?             H@������������������������       �R�}e�.�?             :@������������������������       �                     6@                           �?      �?             0@������������������������       ��θ�?	             *@������������������������       �                     @        #                    @~�EH,��?d            �b@!       "                   �_@��}*_��?7            @T@������������������������       �                     "@������������������������       ��q�q�?2             R@$       %                   `s@ ���g=�?-            @Q@������������������������       ��C��2(�?*            �P@������������������������       ��q�q�?             @'       ,                    �?<���D�?9            �X@(       +                   �r@      �?             6@)       *       	          ���@     ��?             0@������������������������       �                     @������������������������       �X�<ݚ�?             "@������������������������       �                     @-       .                   �r@�e���@�?.            @S@������������������������       �        %             O@/       0                    �O@��S�ۿ?	             .@������������������������       �                     $@������������������������       �z�G�z�?             @�t�bh�h(h+K ��h-��R�(KK1KK��ha�B        q@     Pu@     �T@     `k@      9@      h@      (@     �e@      "@     �e@      "@     �F@              `@      @              *@      3@      @      3@      @                      3@      "@              M@      :@      @@              :@      :@      @      4@      @               @      4@      5@      @      2@              @      @     �g@     �^@      Z@     �[@      *@     �I@      @     �D@      @      3@              6@      @      $@      @      $@      @             �V@     �M@      >@     �I@      "@              5@     �I@     �N@       @      N@      @      �?       @     �U@      (@      &@      &@      @      &@              @      @      @      @              S@      �?      O@              ,@      �?      $@              @      �?�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ���hG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK-hyh(h+K ��h-��R�(KK-��h��B�	                             �?�:�Ӛ��?�           8�@                          �p@�>ټʹ�?�            `s@       
                    �?�
���?r            �g@                           �?N{�T6�?             �K@                           �?�MI8d�?            �B@������������������������       �                     ;@������������������������       ����Q��?             $@       	                    @r�q��?
             2@������������������������       �      �?             @������������������������       �                     (@                           �?��M���?R             a@                           �?�q�����?              I@������������������������       ����y4F�?             3@������������������������       �f���M�?             ?@                           \@�T|n�q�?2            �U@������������������������       �X�<ݚ�?
             2@������������������������       �l��\��?(             Q@                          �b@��u}���?J            �]@                           @ ��N8�?3             U@                          Ps@      �?             @@������������������������       ��C��2(�?
             &@������������������������       �        
             5@������������������������       �                     J@                           �?4�2%ޑ�?            �A@              	          ����?X�<ݚ�?             2@������������������������       ��n_Y�K�?             *@������������������������       �                     @������������������������       �        	             1@       ,                    g@��^͝B�?�            s@       %                    @ ��-{F�?�            �r@       "                    �?T�W2��?�            �m@        !                    �?p�ݯ��?             3@������������������������       �                     (@������������������������       �                     @#       $                   �_@F��}��?�            `k@������������������������       ��q�q�?             (@������������������������       ���+��?�            �i@&       )       	          `ff�?4�.�A�?.            �O@'       (                    @I@      �?"             F@������������������������       �և���X�?             @������������������������       ���G���?            �B@*       +       
             �?���y4F�?             3@������������������������       �                     @������������������������       �        
             .@������������������������       �                     @�t�bh�h(h+K ��h-��R�(KK-KK��ha�B�       `q@     u@     �l@     @T@     �]@      R@      5@      A@      @      ?@              ;@      @      @      .@      @      @      @      (@             �X@      C@      :@      8@      .@      @      &@      4@      R@      ,@      $@       @      O@      @     �[@      "@     �T@      �?      ?@      �?      $@      �?      5@              J@              ;@       @      $@       @      @       @      @              1@             �H@      p@     �F@      p@      3@     `k@      @      (@              (@      @              (@     �i@      @       @       @     �h@      :@     �B@      &@     �@@      @      @      @      >@      .@      @              @      .@              @        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJJ��hG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK3hyh(h+K ��h-��R�(KK3��h��B(                             �?��>�'��?�           8�@                           @d�B��?           0y@       
       	          033�?�A����?�            @q@                          �s@�cX1!��?�             o@                           @L@=QcG��?�            `m@������������������������       ��d���?k            �e@������������������������       �L=�m��?,            �N@       	                    @L@X�Cc�?             ,@������������������������       �                     @������������������������       �X�<ݚ�?             "@                           @F@|��?���?             ;@������������������������       �                     @                          �_@��Q��?             4@������������������������       �r�q��?             @������������������������       �؇���X�?	             ,@                           �?fȮ�Б�?P            �_@              	          ����?�S����?"            �L@                           �O@�q�q�?             ;@������������������������       ���+7��?             7@������������������������       �      �?             @������������������������       �                     >@              	          ����?��(@��?.            �Q@              
             �?0,Tg��?             E@������������������������       ��G�z��?             4@������������������������       ��C��2(�?             6@              	          ���@d}h���?             <@������������������������       �H%u��?             9@������������������������       �                     @       *       	          ����?���U�?�            �j@       %                    @P�=?!�?@            @[@       "                    �?l��[B��?$             M@        !                   �n@�������?             A@������������������������       �      �?              @������������������������       �8�Z$���?             :@#       $                    �?�q�q�?             8@������������������������       �      �?             $@������������������������       �                     ,@&       )       	          pff�?��x_F-�?            �I@'       (                    �?X�Cc�?             <@������������������������       ������H�?             "@������������������������       ��\��N��?
             3@������������������������       �                     7@+       0                    @�]��?F            �Y@,       /                    �F@p���?C             Y@-       .       	          033@�t����?             1@������������������������       �        	             ,@������������������������       ��q�q�?             @������������������������       �        7            �T@1       2                    �I@�q�q�?             @������������������������       �                     �?������������������������       �                      @�t�bh�h(h+K ��h-��R�(KK3KK��ha�B0       �q@     �t@     �\@     r@     �@@     `n@      4@     �l@      .@     �k@      @     @e@      &@      I@      @      "@              @      @      @      *@      ,@              @      *@      @      �?      @      (@       @     @T@      G@      H@      "@      2@      "@      1@      @      �?      @      >@             �@@     �B@      &@      ?@      "@      &@       @      4@      6@      @      6@      @              @     @e@      E@     �Q@      C@      >@      <@      9@      "@      @      @      6@      @      @      3@      @      @              ,@     �D@      $@      2@      $@       @      �?      $@      "@      7@             �X@      @     �X@       @      .@       @      ,@              �?       @     �T@              �?       @      �?                       @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ�U�uhG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK3hyh(h+K ��h-��R�(KK3��h��B(                             �?�:�Ӛ��?y           8�@              
             �?��5Е��?�            �p@                           @n�tv?�?p            �f@              
             �?4�B��?-            �R@������������������������       �                     &@                           b@�ՙ/�?&            �O@������������������������       ���
ц��?             J@������������������������       �                     &@	                           �O@�8�l��?C            �Z@
                          �c@�L��ȕ?;            @W@������������������������       �        5            �T@������������������������       �ףp=
�?             $@                          (p@��
ц��?             *@������������������������       �                     @������������������������       �                     @                           �?X�����?7             V@                          0f@      �?             H@������������������������       �                     @                          �c@"pc�
�?             F@������������������������       �ҳ�wY;�?	             1@������������������������       ��>����?             ;@                           �?z�G�z�?             D@                           �?�q�q�?             5@������������������������       �                     @������������������������       �        	             ,@������������������������       �                     3@       *       	          033�?xO.�|�?�            �u@       #                    @�h�]���?�            pr@               
             �?�K�w���?�            `l@                           �?���N8�?%            �O@������������������������       �@3����?             K@������������������������       ��<ݚ�?             "@!       "                    �?�qE��E�?f            �d@������������������������       ����-T��?'             O@������������������������       ��IєX�??            �Y@$       '                    �?j���� �?*             Q@%       &                   8p@f.i��n�?            �F@������������������������       �ܷ��?��?             =@������������������������       �     ��?	             0@(       )                    �?�û��|�?             7@������������������������       ��q�q�?             5@������������������������       �                      @+       ,                   �[@R�}e�.�?             J@������������������������       �                     @-       0                     G@�㙢�c�?             G@.       /                   �e@z�G�z�?             @������������������������       �                     @������������������������       �                     �?1       2                    b@������?            �D@������������������������       �P�Lt�<�?             C@������������������������       �                     @�t�bh�h(h+K ��h-��R�(KK3KK��ha�B0       `q@     u@     @h@     �R@     �b@      ?@      I@      8@      &@             �C@      8@      <@      8@      &@             �X@      @      W@      �?     �T@              "@      �?      @      @      @                      @     �F@     �E@      (@      B@      @               @      B@      @      &@       @      9@     �@@      @      ,@      @              @      ,@              3@              U@     pp@      G@      o@      2@      j@      @      N@      �?     �J@       @      @      .@     �b@      "@     �J@      @      X@      <@      D@      ,@      ?@      @      :@      &@      @      ,@      "@      ,@      @               @      C@      ,@              @      C@       @      �?      @              @      �?             �B@      @     �B@      �?              @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJW��]hG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK1hyh(h+K ��h-��R�(KK1��h��B�
                             �?�p ��?�           8�@                           �?,N��tf�?�            �x@       
                    �?T���RB�?�             o@                           @ܩ�d	��?,            �S@                          �`@4և����?!             L@������������������������       ��חF�P�?             ?@������������������������       �                     9@       	                    @K@8����?             7@������������������������       ��S����?             3@������������������������       �                     @                          �[@<���i�?j            @e@                          �k@      �?             @@������������������������       �                     ,@������������������������       ��q�q�?	             2@                           @@��9U��?Z            @a@������������������������       ��g�y��?R             _@������������������������       �d}h���?             ,@              	          ����?��ӭ�a�?b             b@                           �?$��m��?6            �S@                          �s@������?            �B@������������������������       ��g�y��?             ?@������������������������       �      �?             @              
             �?�>$�*��?            �D@������������������������       �      �?             (@������������������������       �8^s]e�?             =@                          �l@r�q��?,            �P@������������������������       �                     >@                           �?<ݚ)�?             B@������������������������       �ףp=
�?             4@������������������������       �     ��?             0@       (                    @���GYW�?�            �k@        !                   �]@�E���?=            @X@������������������������       �                     :@"       %                    �?`��_��?,            �Q@#       $                    �?f.i��n�?            �F@������������������������       �      �?
             0@������������������������       �\-��p�?             =@&       '                    �?8�Z$���?             :@������������������������       �        	             ,@������������������������       ��q�q�?             (@)       *                   �Z@H�̱���?N            @_@������������������������       �                     @+       .                   �[@ �p���?L            �^@,       -                    Z@PN��T'�?             ;@������������������������       �                     *@������������������������       �����X�?             ,@/       0                    �?�eGk�T�?:            �W@������������������������       � ��N8�?4             U@������������������������       �                     &@�t�bh�h(h+K ��h-��R�(KK1KK��ha�B       �r@     �s@     �^@     �p@      D@      j@      5@      M@      @     �I@      @      :@              9@      0@      @      0@      @              @      3@     �b@      (@      4@              ,@      (@      @      @     ``@      @      ^@      @      &@     �T@      O@      ;@     �I@      @     �@@      �?      >@      @      @      7@      2@      @      "@      4@      "@     �K@      &@      >@              9@      &@      2@       @      @      "@     @f@      F@     �N@      B@      :@             �A@      B@      ?@      ,@      @      $@      9@      @      @      6@              ,@      @       @     @]@       @              @     @]@      @      7@      @      *@              $@      @     �W@      �?     �T@      �?      &@        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJt�mUhG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK/hyh(h+K ��h-��R�(KK/��h��BH
                             �?;�׊��?}           8�@                           �?�=Aq�4�?�            @s@              	          pff�?>��T��?W            �a@                           �D@h/��y��?-            @S@������������������������       �                     @                          �n@�q�q�?)             R@������������������������       �X�EQ]N�?            �E@������������������������       �J�8���?             =@	                           @��s����?*            �O@
              	          033�?p�ݯ��?             3@������������������������       �8�Z$���?
             *@������������������������       �r�q��?             @������������������������       �                     F@                          �Z@�h����?f             e@                           �?z�G�z�?
             $@                           Y@����X�?             @������������������������       �                     @������������������������       ��q�q�?             @������������������������       �                     @              	          ����?��o;���?\            �c@                           �?8��8���?             H@������������������������       ���a�n`�?             ?@������������������������       �                     1@������������������������       �        @            �[@       (       	          033�?��2p��?�            0s@       !       
             �?V���w�?�            Pq@                          �[@z�G�z�?7            @U@              	          pff�?      �?             $@������������������������       �r�q��?             @������������������������       �                     @                            �K@�J�4�?0            �R@������������������������       ��?�|�?            �B@������������������������       �p9W��S�?             C@"       %                    �?�8��8��?u             h@#       $                   f@����?+            �S@������������������������       �                     @������������������������       �DE��2{�?)            �R@&       '                   c@�}�+r��?J            �\@������������������������       ���<b���?             7@������������������������       �@��,B�?=            �V@)       .                    �?z�G�z�?             >@*       +       	          `ff@���Q��?             $@������������������������       �                     @,       -                   g@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     4@�t�bh�h(h+K ��h-��R�(KK/KK��ha�B�       �r@     �s@     �l@     �S@     �Q@     @Q@      4@     �L@      @              .@     �L@      @      C@      $@      3@     �I@      (@      @      (@       @      &@      @      �?      F@             �c@      "@       @       @      @       @      @              �?       @      @             �b@      @     �D@      @      8@      @      1@             �[@             �P@      n@      E@     `m@      1@      Q@      @      @      @      �?              @      (@     �O@      �?      B@      &@      ;@      9@     �d@      3@     �M@      @              0@     �M@      @      [@      @      2@      �?     �V@      8@      @      @      @              @      @      �?      @                      �?      4@        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJc��hG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK/hyh(h+K ��h-��R�(KK/��h��BH
                             �?��O���?�           8�@                           �?P�r;�?           �y@       
       	          033�?�L����?�            @o@                           @؇���X�?�            �m@                           @M@������?y            @f@������������������������       ��J�T�?]            �a@������������������������       ��E��ӭ�?             B@       	                    �?�q�q�?%             N@������������������������       �                      @������������������������       ��n_Y�K�?"             J@                           �?�q�q�?             (@������������������������       �                     @                           �E@      �?              @������������������������       �                     @������������������������       �      �?             @              
             �?��y���?]            �c@                           @G@ڤ���?.            @T@������������������������       �                     @                          �a@��n�?,            �R@������������������������       �$�q-�?            �C@������������������������       �<ݚ)�?             B@                           f@\I�~�?/            @S@                           �P@      �?-             R@������������������������       ���o	��?&             M@������������������������       �                     ,@������������������������       �                     @       (                    �?�! *��?�            �i@       !                    �?���I�?q            `f@               	          ����?���@��?            �B@              	          ����?�n_Y�K�?             *@������������������������       �      �?              @������������������������       �                     @������������������������       �                     8@"       %                   �Z@,�d�vK�?[            �a@#       $                   �Y@���Q��?             @������������������������       �                      @������������������������       �                     @&       '                   �d@A_�&�?W             a@������������������������       ��wY;��?V             a@������������������������       �                     �?)       *                   �\@X�Cc�?             <@������������������������       �                     @+       .       	             �?�eP*L��?             6@,       -                   0o@$�q-�?
             *@������������������������       �                     &@������������������������       �      �?              @������������������������       �                     "@�t�bh�h(h+K ��h-��R�(KK/KK��ha�B�        s@     ps@     �`@      q@     �D@      j@      A@     �i@      ,@     �d@      @     @a@      $@      :@      4@      D@               @      4@      @@      @      @      @              @      @              @      @      �?     @W@     @P@     �N@      4@              @     �N@      ,@      B@      @      9@      &@      @@     �F@      ;@     �F@      ;@      ?@              ,@      @             @e@     �B@      d@      3@      =@       @      @       @      @      @              @      8@             ``@      &@       @      @       @                      @      `@       @      `@      @              �?      $@      2@              @      $@      (@      �?      (@              &@      �?      �?      "@        �t�bubhhubh)��}�(hhhhhKhKhKhG        �P	     hh$hNhJg�$hG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK3hyh(h+K ��h-��R�(KK3��h��B(                             @f�*�L�?�           8�@              	          033�?�̫+ 4�?�            px@       
                    �?H~4o]�?�            �u@                          Pb@���-|$�?`            @c@                           �?�Ƀ aA�?#            �M@������������������������       ��8��8��?             8@������������������������       �^������?            �A@       	                    a@\�ih�<�?=            �W@������������������������       �d}h���?'             L@������������������������       � ���J��?            �C@                          �d@     �?r             h@                           �? 7���B�?p            �g@������������������������       �pY���D�?[            �c@������������������������       ���a�n`�?             ?@                          �q@�q�q�?             @������������������������       �                      @������������������������       �                     �?                           @O@:	��ʵ�?            �F@                           �?�8��8��?             B@������������������������       �                     2@              
             �?r�q��?             2@������������������������       ��t����?             1@������������������������       �                     �?                           �?X�<ݚ�?             "@������������������������       �                     @                          0a@z�G�z�?             @������������������������       ��q�q�?             @������������������������       �                      @       (       	          pff�?���>4��?�             l@       %                   �p@�Je\���?3            @T@       "                   �^@      �?'             P@        !                    �?؇���X�?             5@������������������������       �                     @������������������������       �z�G�z�?	             .@#       $                    �?X��ʑ��?            �E@������������������������       ��ʻ����?             A@������������������������       ��<ݚ�?             "@&       '                   �a@�IєX�?             1@������������������������       �                     �?������������������������       �                     0@)       .       	          ����?�C����?a            �a@*       -                   X{@�Q��k�?5             T@+       ,                   pb@��r�Z}�?4            �S@������������������������       �lGts��?%            �K@������������������������       �      �?             8@������������������������       �                     �?/       0                    @M@ ������?,            �O@������������������������       �                    �B@1       2                   �p@ ��WV�?             :@������������������������       �                     4@������������������������       �r�q��?             @�t�bh�h(h+K ��h-��R�(KK3KK��ha�B0       `p@     v@     @W@     �r@      L@      r@     �G@     �Z@      A@      9@      6@       @      (@      7@      *@     �T@      (@      F@      �?      C@      "@     �f@      @     �f@      @     @c@      @      <@       @      �?       @                      �?     �B@       @     �@@      @      2@              .@      @      .@       @              �?      @      @              @      @      �?       @      �?       @              e@     �K@      D@     �D@      8@      D@      @      2@              @      @      (@      5@      6@      3@      .@       @      @      0@      �?              �?      0@              `@      ,@     �P@      *@     �P@      (@     �H@      @      2@      @              �?      O@      �?     �B@              9@      �?      4@              @      �?�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ�>D5hG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK3hyh(h+K ��h-��R�(KK3��h��B(                
             �?���>��?�           8�@                          pb@�^�����?�            �u@       
                    �?lkч��?�            �m@                           �?0d4�[%�?;            �W@                           �P@D�n�3�?             C@������������������������       ��g�y��?             ?@������������������������       �                     @       	                   i@���5��?#            �L@������������������������       �                     :@������������������������       ���a�n`�?             ?@                           �?�X�<ݺ?Q             b@������������������������       �        1            �U@              	          ����?Ԫ2��?             �L@������������������������       �                     @������������������������       �`'�J�?            �I@              	          pff�?n�����?D            @Z@                           @ȵHPS!�?"             J@������������������������       �                     C@                          @d@և���X�?	             ,@������������������������       ����!pc�?             &@������������������������       �                     @                           @Fmq��?"            �J@              	          `ff
@      �?             8@������������������������       �؇���X�?             5@������������������������       �                     @                          X~@ܷ��?��?             =@������������������������       � 7���B�?             ;@������������������������       �                      @       (                    @L@��Vu���?�            �p@       #                    �?4��?�?h            �c@       "                   8q@�%^�?            �E@        !                    �?:�&���?            �C@������������������������       ������H�?             B@������������������������       �                     @������������������������       �                     @$       '                   c@�/�z{�?N            @\@%       &                   �d@�	j*D�?
             *@������������������������       �                      @������������������������       �"pc�
�?	             &@������������������������       �        D             Y@)       .                    @~}e}b �?H            �\@*       -                   @e@����X�?/            @S@+       ,                    �?��>4և�?$             L@������������������������       �j���� �?             A@������������������������       ��C��2(�?             6@������������������������       �                     5@/       0                    �?�����?             C@������������������������       �                      @1       2                     P@�E��ӭ�?             B@������������������������       ��חF�P�?             ?@������������������������       �                     @�t�bh�h(h+K ��h-��R�(KK3KK��ha�B0       �r@     �s@      n@      Z@     @i@     �B@     �P@      =@      0@      6@      0@      .@              @      I@      @      :@              8@      @      a@       @     �U@             �H@       @              @     �H@       @      C@     �P@      @      G@              C@      @       @      @       @      @              @@      5@      @      2@      @      2@      @              :@      @      :@      �?               @     �O@      j@      .@     �a@      &@      @@      @      @@      @      @@      @              @              @     @[@      @      "@       @               @      "@              Y@      H@     �P@      6@     �K@      6@      A@      4@      ,@       @      4@              5@      :@      (@               @      :@      $@      :@      @              @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ���&hG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK/hyh(h+K ��h-��R�(KK/��h��BH
                	          033�?��>�'��?�           8�@                           @8�zJ�?&            }@       
                    �?BK"(<\�?�            0t@                          �`@ҳ�wY;�?G            �]@                          `f@$/����?,            @P@������������������������       �П[;U��?'             M@������������������������       �                     @       	                   0b@�+$�jP�?             K@������������������������       �                     $@������������������������       �                     F@                          �d@l��\��?�            �i@                           �?Riv����?K             ]@������������������������       ��~i��?E            @[@������������������������       �؇���X�?             @������������������������       �        9             V@                           �?"Ae���?[            �a@                          @[@��2(&�?8             V@                           Z@      �?             @������������������������       �                     �?������������������������       �                     @              	          ����? �Cc}�?6             U@������������������������       �      �?             B@������������������������       �                     H@                          �b@`��}3��?#            �J@              	          833�?�eP*L��?             6@������������������������       ��θ�?             *@������������������������       �                     "@                           �?�חF�P�?             ?@������������������������       �      �?             $@������������������������       �                     5@       $                    �F@�ș�j�?[            �b@        #                    @8�A�0��?             6@!       "                    �?X�Cc�?             ,@������������������������       �                     @������������������������       �                     "@������������������������       �                      @%       *                    �?,mG����?N             `@&       )                    @�㙢�c�?              G@'       (                    �?�����?             E@������������������������       �h�����?             <@������������������������       �d}h���?             ,@������������������������       �                     @+       ,                    �O@P��BNֱ?.            �T@������������������������       �        %             P@-       .                    �?�S����?	             3@������������������������       ����Q��?             @������������������������       �                     ,@�t�bh�h(h+K ��h-��R�(KK/KK��ha�B�       �q@     �t@      c@     ps@      N@     pp@      E@     @S@      @@     �@@      @@      :@              @      $@      F@      $@                      F@      2@     @g@      2@     �X@      (@     @X@      @      �?              V@     @W@      H@      S@      (@      �?      @      �?                      @     �R@      "@      ;@      "@      H@              1@      B@      (@      $@      @      $@      "@              @      :@      @      @              5@     ``@      4@      *@      "@      @      "@      @                      "@       @             �]@      &@      C@       @      C@      @      ;@      �?      &@      @              @      T@      @      P@              0@      @       @      @      ,@        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ�EhG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK7hyh(h+K ��h-��R�(KK7��h��B                             �?Z�����?�           8�@              
             �?��t�%�?�            ps@       
                   pb@r�q��?�            @j@                           �?��㨇,�?i            �e@                           �?��<b�ƥ?8             W@������������������������       �r�q��?             (@������������������������       �        0             T@       	       	          ����?�<ݚ�?1            @T@������������������������       ��q�q�?             .@������������������������       �<���D�?)            �P@              	             �?�Gi����?            �B@                           �?8�Z$���?	             *@������������������������       ��8��8��?             (@������������������������       �                     �?                          �e@r�q��?             8@������������������������       ��C��2(�?             6@������������������������       �                      @                          0f@:�o���?7            @Y@                           @ 9�����?1             V@                           �?p�v>��?            �G@������������������������       �                     @������������������������       ��X����?             F@                           �?� ��1�?            �D@������������������������       ��q�q�?	             (@������������������������       �XB���?             =@������������������������       �                     *@       (                   �a@���y4F�?�             s@       #                    �?X�Emq�?#            �J@                           �_@���!pc�?             6@                           @z�G�z�?             @������������������������       �                     �?������������������������       �                     @!       "                   `c@�t����?             1@������������������������       �                     .@������������������������       �                      @$       %       	          ����?��a�n`�?             ?@������������������������       �                     @&       '                   hr@؇���X�?             <@������������������������       �`2U0*��?             9@������������������������       �                     @)       0                   c@@�g8���?�            `o@*       -                    �? �o_��?!             I@+       ,                    �?�������?             F@������������������������       �        	             1@������������������������       ��q�q�?             ;@.       /                    �?r�q��?             @������������������������       �      �?              @������������������������       �                     @1       4                    �?����#��?�             i@2       3       
             �?@	tbA@�?/            @Q@������������������������       �P���Q�?             4@������������������������       �                     �H@5       6                   ``@�禺f��?U            �`@������������������������       ��X�<ݺ?2             R@������������������������       �      �?#             N@�t�bh�h(h+K ��h-��R�(KK7KK��ha�Bp       �q@     �t@     �k@     @V@     �e@     �A@      c@      4@     �V@       @      $@       @      T@             �O@      2@      @      $@      M@       @      6@      .@       @      &@      �?      &@      �?              4@      @      4@       @               @     �G@      K@     �G@     �D@      ,@     �@@              @      ,@      >@     �@@       @      @      @      <@      �?              *@      P@      n@      >@      7@      @      0@      @      �?              �?      @               @      .@              .@       @              8@      @              @      8@      @      8@      �?              @      A@      k@      ,@      B@      "@     �A@              1@      "@      2@      @      �?      �?      �?      @              4@     �f@      �?      Q@      �?      3@             �H@      3@     @\@      @      Q@      .@     �F@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ4�phG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK3hyh(h+K ��h-��R�(KK3��h��B(                             �?*�3�V��?v           8�@                           �?��x/4��?�            0z@       
       	          ����?tv?z���?k            �f@                           �?��x�5��?X            @a@                          `f@�Q��k�?/             T@������������������������       �                     @������������������������       ���}���?-            @S@       	                    w@�BbΊ�?)             M@������������������������       �D>�Q�?&             J@������������������������       �                     @                           @�����?             E@                           �? ���J��?            �C@������������������������       �                     �?������������������������       �                     C@������������������������       �                     @              	          033�?P��8�?�            �m@                           @�W��?�            �k@                          @[@�8��8��?`             e@������������������������       ��<ݚ�?
             2@������������������������       ���S�ۿ?V            �b@              	          ����?`��}3��?$            �J@������������������������       �tk~X��?             B@������������������������       �j���� �?             1@              
             �?�����H�?             2@                           q@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �        
             .@       &       	          ����?Jm_!'1�?{            �h@       %                    �?
;&����?             G@       "       
             �?��Zy�?            �C@        !                    p@�t����?	             1@������������������������       �                     (@������������������������       �                     @#       $                   `d@�GN�z�?             6@������������������������       �     ��?
             0@������������������������       �                     @������������������������       �                     @'       .                    �?���Lͩ�?_            �b@(       +       	          pff�?��J��i�?U            �`@)       *                   �s@�q�q�?             @������������������������       �                      @������������������������       �                     �?,       -                   �j@@��A1ʞ?R            ``@������������������������       �@9G��?            �H@������������������������       �        6            �T@/       0       	          ����?     ��?
             0@������������������������       �                      @1       2                    �?d}h���?	             ,@������������������������       �                     @������������������������       ����!pc�?             &@�t�bh�h(h+K ��h-��R�(KK3KK��ha�B0       �r@     �s@     �a@     `q@     �W@     �U@      L@     �T@      *@     �P@      @              $@     �P@     �E@      .@     �E@      "@              @      C@      @      C@      �?              �?      C@                      @     �G@      h@      ?@     �g@      ,@     @c@      @      ,@      $@     �a@      1@      B@      @      =@      $@      @      0@       @      �?       @               @      �?              .@              d@      B@      8@      6@      1@      6@      (@      @      (@                      @      @      1@      @      &@              @      @              a@      ,@     ``@      @       @      �?       @                      �?      `@       @     �G@       @     �T@              @      &@       @              @      &@              @      @       @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJLxhG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK7hyh(h+K ��h-��R�(KK7��h��B                             �?b�#�(��?�           8�@              	          pff�?�%t�l-�?�            �p@       
                    @���ջ��?E             Z@                           �?�z�G��?*             N@                            N@ףp=
�?             D@������������������������       �                     >@������������������������       ����Q��?             $@       	                    �?�z�G��?             4@������������������������       ��<ݚ�?             2@������������������������       �                      @                          �^@v�X��?             F@                           Z@�<ݚ�?             "@������������������������       �                     �?������������������������       �      �?              @                           @O@b�h�d.�?            �A@������������������������       ���a�n`�?             ?@������������������������       �      �?             @                           �?��1���?m            �d@������������������������       �        =            �T@                           f@R�(CW�?0            �T@                          0s@ȵHPS!�?-            �S@������������������������       �@�r-��?#            �M@������������������������       �        
             3@������������������������       �                     @       (       
             �?"��Ƥ��?�            �u@       !                    �K@�Z4���?M            �`@                           @h��Q(�?'            �P@                          @^@���5��?             �L@������������������������       �H�V�e��?             A@������������������������       �                     7@                            @H@�z�G��?             $@������������������������       �                     @������������������������       �                     @"       %                    �?���`��?&            �P@#       $       
             �?4�B��?            �B@������������������������       �                     "@������������������������       �և���X�?             <@&       '                   �a@z�G�z�?             >@������������������������       �д>��C�?             =@������������������������       �                     �?)       0                   c@�����?�            �j@*       -                    �?������?              L@+       ,                   @[@؇���X�?             E@������������������������       �                      @������������������������       �ףp=
�?             D@.       /                    �?@4և���?             ,@������������������������       �                     *@������������������������       �                     �?1       4                   �t@��)�G��?e            �c@2       3       	          hff@�w�uz
�?^            �a@������������������������       �`�q�0ܴ?\            �a@������������������������       �                      @5       6                    �?�θ�?             *@������������������������       ����!pc�?             &@������������������������       �                      @�t�bh�h(h+K ��h-��R�(KK7KK��ha�Bp       �q@     �t@      i@      Q@     �H@     �K@      2@      E@      @      B@              >@      @      @      ,@      @      ,@      @               @      ?@      *@       @      @      �?              �?      @      =@      @      <@      @      �?      @      c@      *@     �T@             @Q@      *@     @Q@      "@      I@      "@      3@                      @      T@     �p@      I@      U@      ,@     �J@      @      I@      @      ;@              7@      @      @      @                      @      B@      ?@      (@      9@              "@      (@      0@      8@      @      8@      @              �?      >@     �f@      3@     �B@      @      B@       @              @      B@      *@      �?      *@                      �?      &@      b@       @     �`@      @     �`@       @              @      $@      @       @               @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJW��8hG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK3hyh(h+K ��h-��R�(KK3��h��B(                            Pb@�85�r��?}           8�@              
             �?�(�Tw��?�            q@                           �?�{��?��?             k@              	          ����?��j��?+            @S@������������������������       �        
             2@                          @\@6�iL�?!            �M@������������������������       �                     @������������������������       ��rF���?            �K@	              	          ����?���۟�?T            `a@
                           `@@�r-��?"            �M@������������������������       ����Q��?             4@������������������������       � ���J��?            �C@                           @@�z�G�?2             T@������������������������       �        1            �S@������������������������       �                     �?                           @D�n�3�?"            �L@                           �K@�w��#��?             I@������������������������       �        	             .@                          �^@��
P��?            �A@������������������������       ��θ�?	             *@������������������������       ����|���?             6@������������������������       �                     @       $                    @Xb>��?�            `u@                          0e@�uD����?�             m@              
             �?V��~��?a            �b@              	          033�?�D��?             �H@������������������������       �                    �A@������������������������       �@4և���?
             ,@                          �s@.p����?A            @Y@������������������������       �xP�Fֺ�?8            @V@������������������������       ��q�q�?	             (@        !                    �?P��BNֱ?7            �T@������������������������       �        ,             P@"       #                    �?�S����?             3@������������������������       �      �?              @������������������������       �                     &@%       ,                    �?�q�QQ�?D            @[@&       )                   `\@f>�cQ�?%            �N@'       (                    �K@��
ц��?             *@������������������������       �      �?              @������������������������       �                     @*       +                   �n@      �?             H@������������������������       �R���Q�?
             4@������������������������       �                     <@-       0                    �?     ��?             H@.       /       	          hff @4���C�?            �@@������������������������       ���X��?             <@������������������������       �                     @1       2                    �?��S�ۿ?             .@������������������������       �$�q-�?             *@������������������������       �                      @�t�bh�h(h+K ��h-��R�(KK3KK��ha�B0       �r@     �s@     �h@     @S@     �e@      F@     �E@      A@              2@     �E@      0@              @     �E@      (@      `@      $@      I@      "@      (@       @      C@      �?     �S@      �?     �S@                      �?      8@     �@@      1@     �@@              .@      1@      2@      @      $@      ,@       @      @             @Y@      n@      A@     �h@      ?@     �]@      *@      B@             �A@      *@      �?      2@     �T@      &@     �S@      @      @      @      T@              P@      @      0@      @      @              &@     �P@      E@      J@      "@      @      @       @      @      @             �F@      @      1@      @      <@              .@     �@@      ,@      3@      "@      3@      @              �?      ,@      �?      (@               @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ��UhG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK1hyh(h+K ��h-��R�(KK1��h��B�
                
             �?�:�Ӛ��?�           8�@                           �?��ҧ��?�            �t@       
                   �e@֦�r���?p            �e@                           �?�j����?g            �c@                          �d@     ��?<             X@������������������������       �U7W1�?5            �T@������������������������       ��	j*D�?             *@       	                    �?X��Oԣ�?+             O@������������������������       ��?�|�?            �B@������������������������       ��+e�X�?             9@������������������������       �        	             ,@                           �?��-�=��?g            �c@                          �Z@HX���?U            ``@                           �M@r�q��?             @������������������������       �                     @������������������������       �                     �?                          �a@HP�s��?R            @_@������������������������       � f^8���?C            �Y@������������������������       ��X����?             6@              	          ����?`2U0*��?             9@                          �a@�����H�?             "@������������������������       �                     @������������������������       ��q�q�?             @������������������������       �                     0@       $                    @L@"&��E�?�            �q@                           @�:�^���?j            �c@                           �?���}��?X            �`@������������������������       �        B            �X@                           �?������?             A@������������������������       �                     @������������������������       � 7���B�?             ;@        !                   g@��+7��?             7@������������������������       �                      @"       #                    �?��s����?             5@������������������������       �      �?             @������������������������       ��IєX�?             1@%       *                   �a@��w��?N            ``@&       '                    �N@� �	��?             9@������������������������       �                     $@(       )                    �?������?             .@������������������������       �                     @������������������������       �X�<ݚ�?             "@+       .                    �?v�XԖ�??            �Z@,       -                   d@      �?             B@������������������������       �      �?             0@������������������������       ��z�G��?             4@/       0                    �?ףp=
�?&            �Q@������������������������       �r�q��?             >@������������������������       �P���Q�?             D@�t�bh�h(h+K ��h-��R�(KK1KK��ha�B       `q@     u@      l@     �Y@     @U@     �U@     @U@     @R@      >@     �P@      5@      O@      "@      @     �K@      @      B@      �?      3@      @              ,@     �a@      0@      ]@      .@      �?      @              @      �?             �\@      $@      Y@      @      .@      @      8@      �?       @      �?      @               @      �?      0@             �J@     @m@      ,@     �a@       @     @_@             �X@       @      :@      @              �?      :@      @      1@       @              @      1@      @      �?      �?      0@     �C@      W@      ,@      &@      $@              @      &@              @      @      @      9@     @T@      2@      2@      @      (@      ,@      @      @     �O@      @      9@       @      C@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ��DphG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK5hyh(h+K ��h-��R�(KK5��h��B�                             �?V���Ş�?�           8�@                           �?�3��f�?�             s@       
                    @���>4��?/             U@                          `a@X�Cc�?%            �Q@              	          ����?�<ݚ�?             K@������������������������       ����Q��?             >@������������������������       �                     8@       	                   �b@     ��?
             0@������������������������       �                     $@������������������������       �      �?             @������������������������       �        
             ,@                           �?���GYW�?�            �k@                           @t�C�#��?8            �S@                           �P@�e����?            �C@������������������������       ��!���?             A@������������������������       �                     @                            P@R���Q�?             D@������������������������       ��C��2(�?            �@@������������������������       �և���X�?             @                          �d@�1�hP	�?U            �a@                          �[@Tۢ��(�?R            �`@������������������������       ��I�w�"�?             C@������������������������       �`�E���?@            @X@                           a@      �?              @������������������������       �                     @������������������������       �                     @       (                    @tt���A�?�            Ps@       #       	          hff @p�U�ʻ�?�            �m@                           �a@�FVQ&�?�            �l@                           �?���y4F�?             C@������������������������       �                     2@������������������������       ����Q��?             4@!       "                   �d@@�.L3خ?{             h@������������������������       ����1j	�?:            �U@������������������������       ����1��?A            �Z@$       '                    @      �?              @%       &                   n@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @)       .       	          ����?�xGZ���?0            �Q@*       -                    �?     ��?             @@+       ,       	          ����?�X����?             6@������������������������       �                     @������������������������       ���S���?             .@������������������������       �                     $@/       2       
             �?>A�F<�?             C@0       1       	          ���@��a�n`�?             ?@������������������������       �XB���?             =@������������������������       �                      @3       4                   �l@և���X�?             @������������������������       �      �?             @������������������������       �                     @�t�bh�h(h+K ��h-��R�(KK5KK��ha�BP        q@     Pu@      k@     @V@     �C@     �F@      9@     �F@      (@      E@      (@      2@              8@      *@      @      $@              @      @      ,@             @f@      F@      I@      =@      0@      7@      &@      7@      @              A@      @      >@      @      @      @      `@      .@      _@      &@      =@      "@     �W@       @      @      @              @      @             �L@     �o@      3@     �k@      ,@      k@       @      >@              2@       @      (@      @     `g@      @     @T@      �?     �Z@      @      @      @      �?      @                      �?               @      C@      @@      @      9@      @      .@              @      @       @              $@      ?@      @      <@      @      <@      �?               @      @      @      @      �?              @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ%�[6hG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK/hyh(h+K ��h-��R�(KK/��h��BH
                             �?�:�Ӛ��?�           8�@              	          033�?��t|�
�?�            y@       
                    @&^�)b�?�            �u@                           @L@     p�?�             p@                           �?@]����?i            @f@������������������������       �        8            �Y@������������������������       �`-�I�w�?1             S@       	                    �?���B���?3            �S@������������������������       ��t����?            �I@������������������������       ��q�q�?             ;@                           �?      �?>             V@                          s@����X�?(             L@������������������������       �������?'             K@������������������������       �                      @                           �I@      �?             @@������������������������       ����Q��?             @������������������������       ��>����?             ;@                          `c@P̏����?$            �L@                          �j@ZՏ�m|�?            �H@������������������������       �                     (@                           �F@���@��?            �B@������������������������       �                     @������������������������       �<���D�?            �@@                           �?      �?              @������������������������       �                      @������������������������       �                     @       (       	          ����?�8l�9��?�            �j@       #                    �?d}h��?F             \@                           �p@\��<�|�?:            �W@                           �?���|���?"            �K@������������������������       ��[�IJ�?            �G@������������������������       �                      @!       "                   Pd@��(\���?             D@������������������������       �P�Lt�<�?             C@������������������������       �                      @$       '                   ``@�IєX�?             1@%       &                    �?r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     &@)       *                   �a@`'�J�?E            �Y@������������������������       �        4            @S@+       .                   �\@�J�4�?             9@,       -                   @[@�q�q�?             @������������������������       ��q�q�?             @������������������������       �                     @������������������������       �                     3@�t�bh�h(h+K ��h-��R�(KK/KK��ha�B�       `q@     u@     �Z@     `r@      P@     �q@      4@     �m@      @     �e@             �Y@      @     �Q@      .@     �O@      @     �F@      "@      2@      F@      F@      D@      0@      D@      ,@               @      @      <@       @      @       @      9@     �E@      ,@     �D@       @      (@              =@       @              @      =@      @       @      @       @                      @     `e@     �E@     @R@     �C@      R@      7@     �A@      4@      ;@      4@       @             �B@      @     �B@      �?               @      �?      0@      �?      @              @      �?                      &@     �X@      @     @S@              5@      @       @      @       @      �?              @      3@        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ�	3 hG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK5hyh(h+K ��h-��R�(KK5��h��B�                             �?JGC8{��?�           8�@              	          033�?������?�            �v@       
                    �?�����?�            �r@                           �?�]?ow�?�            �n@                           �?���L��?;            �V@������������������������       �      �?             8@������������������������       �        -            �P@       	                   0b@0z���?`             c@������������������������       ��X����?             6@������������������������       ���ϻ�r�?Q            ``@                          �b@�F�j��?#            �J@                          @]@r֛w���?             ?@������������������������       �                     @������������������������       ��>4և��?             <@                           `@"pc�
�?             6@������������������������       ��q�q�?             "@������������������������       �$�q-�?	             *@                           @M@     ��?$             P@                          �j@ȵHPS!�?             J@                           �?��+7��?             7@������������������������       ���
ц��?             *@������������������������       �                     $@������������������������       �                     =@                          �b@      �?	             (@                           �?�q�q�?             "@������������������������       �                     @������������������������       �                     @������������������������       �                     @       (       	          033�?����H�?�            �o@       #                    �?��F�j�?C            �Z@       "                   @`@�	j*D�?            �C@        !                   �_@X�<ݚ�?             ;@������������������������       �������?             1@������������������������       �z�G�z�?             $@������������������������       �                     (@$       %                    �?D|U��@�?)            �P@������������������������       �                      @&       '                   `g@�?�<��?(            @P@������������������������       �     ��?'             P@������������������������       �                     �?)       .                    �?|��+�?[            �b@*       -                    @�?�|�?D            �[@+       ,                    �?��p\�?            �D@������������������������       �                    �A@������������������������       �      �?             @������������������������       �        +            �Q@/       2                   �l@��+��?            �B@0       1                    �?@4և���?	             ,@������������������������       �                     *@������������������������       �                     �?3       4                   �p@��+7��?             7@������������������������       ����Q��?             .@������������������������       �                      @�t�bh�h(h+K ��h-��R�(KK5KK��ha�BP       �q@     �t@      ]@     �n@      P@      m@     �B@     �i@      @     @U@      @      2@             �P@      ?@     �^@      .@      @      0@     �\@      ;@      :@      7@       @              @      7@      @      @      2@      @      @      �?      (@      J@      (@      G@      @      1@      @      @      @      $@              =@              @      @      @      @              @      @              @             �d@     �V@     �B@     @Q@      ;@      (@      .@      (@      *@      @       @       @      (@              $@     �L@       @               @     �L@      @     �L@      �?             �_@      5@      [@      @      C@      @     �A@              @      @     �Q@              3@      2@      *@      �?      *@                      �?      @      1@      @      "@               @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ��.hG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK3hyh(h+K ��h-��R�(KK3��h��B(                             @Pf�.���?�           8�@                           �J@n^�AL�?�            �w@                           �?���Cu��?j            �d@������������������������       �        +            �Q@                           �?�Ι����??            @X@                           �?�q�q�?             (@������������������������       �                     @������������������������       ��q�q�?             @	       
                    �?�t����?:            @U@������������������������       �      �?             @@������������������������       ��&=�w��?%            �J@                           �?��+�r��?�            �j@                           �?����?8            @V@                           �?     ��?             @@������������������������       �z�G�z�?             4@������������������������       ��8��8��?             (@                          @b@P̏����?#            �L@������������������������       �@4և���?             E@������������������������       �������?
             .@              	              @���N8�?L            �_@                           �M@p�̔B��?D            @\@������������������������       �     ��?%             P@������������������������       �@�E�x�?            �H@                          �a@8�Z$���?             *@������������������������       �                     &@������������������������       �                      @       *       	          ����?��D�^��?�             m@       #                   pc@Rg��J��?@            �X@                            �?�LQ�1	�?             G@                          Pq@z�G�z�?             @������������������������       �                     @������������������������       �                     �?!       "                    �?������?            �D@������������������������       ���.k���?             1@������������������������       �r�q��?             8@$       '                    �?�	j*D�?$             J@%       &                    g@�������?             F@������������������������       ��θ�?            �C@������������������������       �                     @(       )                   �^@      �?              @������������������������       �                     @������������������������       �      �?             @+       ,                    �?�r����?\            �`@������������������������       �                     2@-       0                   �b@8�Z$���?O            @]@.       /                   �e@����"$�?<            �U@������������������������       ���`qM|�?;            �T@������������������������       �                     @1       2                   �a@f���M�?             ?@������������������������       �                     0@������������������������       �������?             .@�t�bh�h(h+K ��h-��R�(KK3KK��ha�B0       �p@     �u@     �Y@     �q@      ,@      c@             �Q@      ,@     �T@      @       @              @      @       @      $@     �R@       @      8@       @     �I@      V@     �_@      M@      ?@      .@      1@      @      0@      &@      �?     �E@      ,@     �C@      @      @      &@      >@      X@      3@     �W@      2@      G@      �?      H@      &@       @      &@                       @      e@      P@      J@      G@      0@      >@      @      �?      @                      �?      (@      =@       @      "@      @      4@      B@      0@     �A@      "@      >@      "@      @              �?      @              @      �?      @     @]@      2@      2@             �X@      2@     �S@      @     �S@      @              @      4@      &@      0@              @      &@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ��~hG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK1hyh(h+K ��h-��R�(KK1��h��B�
                             �?BM�e�x�?           8�@                           �?��B�'m�?�            w@       
                    @L@�wz�~�?�            �q@                           �?��'cy�?y            @i@                          0b@     ��?*             P@������������������������       �      �?             @������������������������       ��8���?$             M@       	                    @@	tbA@�?O            @a@������������������������       �        C            �\@������������������������       ��8��8��?             8@              	          pff�?��X��?2             U@                          �^@     ��?             @@������������������������       �                     @������������������������       ���}*_��?             ;@                          0c@���B���?             J@������������������������       ��t����?             A@������������������������       �        
             2@                          `b@=&C��?3            �T@                           �G@f1r��g�?            �J@������������������������       �                     4@                           �?r٣����?            �@@������������������������       �V�a�� �?             =@������������������������       �      �?             @                           �?�z�G��?             >@������������������������       �                     &@                           @�\��N��?             3@������������������������       �                     @������������������������       �      �?             (@       (                    �?@����]�?�            �n@       #       
             �? 	��p�?d             b@       "                    `@�94�s0�?L            �\@        !                   �_@�:�^���?            �F@������������������������       �                    �B@������������������������       �      �?              @������������������������       �        .            �Q@$       '                   �c@z�G�z�?             >@%       &                    �?և���X�?             ,@������������������������       �      �?              @������������������������       �                     @������������������������       �                     0@)       0       	          033�?�7�yHx�?=            @Y@*       -                   xq@�+e�X�?0            �R@+       ,                    �?PN��T'�?$             K@������������������������       �X�<ݚ�?             2@������������������������       �                     B@.       /                   Hr@�G��l��?             5@������������������������       �                     @������������������������       �������?             .@������������������������       �                     :@�t�bh�h(h+K ��h-��R�(KK1KK��ha�B       �p@     �u@     @V@     �q@     �A@     `o@       @     @h@      @      M@      @      @      @     �K@       @      a@             �\@       @      6@      ;@     �L@      1@      .@              @      1@      $@      $@      E@      $@      8@              2@      K@      =@     �F@       @      4@              9@       @      7@      @       @       @      "@      5@              &@      "@      $@              @      "@      @     `f@     �P@     �`@      $@     �[@      @     �D@      @     �B@              @      @     �Q@              8@      @       @      @       @      @      @              0@              F@     �L@      2@     �L@       @      G@       @      $@              B@      $@      &@      @              @      &@      :@        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ��.hG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK5hyh(h+K ��h-��R�(KK5��h��B�                
             �?��S���?�           8�@                           �?���&#�?�            �t@       
                    @L@`��b���?k            `c@              	          ����?؇>���?/            @P@                           �?@4և���?             E@������������������������       ��q�q�?             @������������������������       �������?             B@       	                    @\X��t�?             7@������������������������       �ףp=
�?             $@������������������������       �$�q-�?             *@              	          pff�?�z�G��?<            �V@                           �P@      �?             8@������������������������       ����y4F�?             3@������������������������       �                     @              
             �?"pc�
�?,            �P@������������������������       ��n_Y�K�?             *@������������������������       �^�!~X�?$            �J@                           �?"pc�
�?l             f@                          �Z@�1�hP	�?Y            �a@              	          033�?      �?             @������������������������       �                     �?������������������������       �                     @                           @��˥W1�?V            `a@������������������������       �     ��?             H@������������������������       �x��B�R�?7            �V@                           �?�'�=z��?            �@@                          �`@`�Q��?             9@������������������������       �                     @������������������������       ��GN�z�?             6@������������������������       �                      @       (                    �?\�CX�?�            �q@        '                   0f@�G�z��?5             T@!       $                    @b�2�tk�?.             R@"       #                   �d@��J�fj�?            �B@������������������������       �������?             ;@������������������������       �ףp=
�?             $@%       &                    @z�G�z�?            �A@������������������������       �6YE�t�?            �@@������������������������       �                      @������������������������       �                      @)       0                    @`�H�/��?�            �i@*       -                   c@��8=��?q            �d@+       ,                    �?z�G�z�?             D@������������������������       �և���X�?             @������������������������       �<���D�?            �@@.       /                    �?`o��b�?U             _@������������������������       � �Jj�G�?&            �K@������������������������       �        /            @Q@1       4                    �?��Q���?             D@2       3                    �?��>4և�?             <@������������������������       ���s����?             5@������������������������       �                     @������������������������       �                     (@�t�bh�h(h+K ��h-��R�(KK5KK��ha�BP       �q@     �t@     �k@      [@     �S@      S@      0@     �H@      @     �C@       @      @      �?     �A@      *@      $@      �?      "@      (@      �?     �O@      ;@      "@      .@      @      .@      @              K@      (@       @      @      G@      @      b@      @@      `@      .@      �?      @      �?                      @     �_@      (@     �C@      "@      V@      @      0@      1@       @      1@      @              @      1@       @              P@     �k@      F@      B@      F@      <@      0@      5@      @      4@      "@      �?      <@      @      <@      @               @               @      4@      g@      "@     `c@       @      @@      @      @      @      =@      �?     �^@      �?      K@             @Q@      &@      =@      &@      1@      @      1@      @                      (@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ�DhG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK7hyh(h+K ��h-��R�(KK7��h��B                
             �?ד�w��?�           8�@                           @R���	�?�             t@       
                    �?���i���?]             c@                           �?����5�?%            �N@                           �?��[�8��?             �I@������������������������       �      �?             6@������������������������       �                     =@       	                    �O@ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?                           �?�y�ʍ+�?8             W@                          `_@     ��?             H@������������������������       �                     @������������������������       �������?            �F@                           �?���7�?             F@������������������������       �؇���X�?	             ,@������������������������       �                     >@                           �?�6���$�?f            �d@              	          ����?      �?0             T@                           `P@8����?             7@������������������������       ����N8�?             5@������������������������       �                      @                           �?l�b�G��?             �L@������������������������       �����X�?             ,@������������������������       �                    �E@                           �O@���E�?6            �U@������������������������       �        ,             S@                           [@�C��2(�?
             &@������������������������       �                     �?������������������������       �        	             $@       ,                   �d@�j;��w�?�            pr@        %                    �?�i�lk��?g            �d@!       "                   �s@�8���?#             M@������������������������       �                    �F@#       $                    �?�θ�?             *@������������������������       �                     $@������������������������       �                     @&       )                    �?����d�?D            @[@'       (                    n@��a�n`�?$             O@������������������������       �      �?             @@������������������������       �*;L]n�?             >@*       +       	          ����?p�v>��?             �G@������������������������       ��}�+r��?             3@������������������������       ����>4��?             <@-       2                   �q@     |�?Y             `@.       1       	          833@@4և���?E            �X@/       0                    �?p�qG�?C             X@������������������������       ��t����?             1@������������������������       �        5            �S@������������������������       �                      @3       4                    �?�q�q�?             >@������������������������       �                     "@5       6                   �d@���N8�?             5@������������������������       �                     4@������������������������       �                     �?�t�bh�h(h+K ��h-��R�(KK7KK��ha�Bp        r@     Pt@     �k@     @X@     @S@      S@      4@     �D@      &@      D@      &@      &@              =@      "@      �?      "@                      �?     �L@     �A@      .@     �@@      @              (@     �@@      E@       @      (@       @      >@             @b@      5@      N@      4@      @      0@      @      0@       @             �J@      @      $@      @     �E@             �U@      �?      S@              $@      �?              �?      $@             �P@     �l@      I@     @]@      @     �K@             �F@      @      $@              $@      @             �G@      O@      ,@      H@      �?      ?@      *@      1@     �@@      ,@      2@      �?      .@      *@      1@     �[@      @     �V@      @     �V@      @      (@             �S@       @              $@      4@      "@              �?      4@              4@      �?        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ���MhG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK=hyh(h+K ��h-��R�(KK=��h��BX                
             �?r � 	��?�           8�@              	          033�?�I� �?�             t@       
                    �?�I{A�?C            �X@                           @؇���X�?*            �O@                           �?ȵHPS!�?"             J@������������������������       ��X�<ݺ?             B@������������������������       �      �?
             0@       	                    �K@���!pc�?             &@������������������������       �                     @������������������������       �և���X�?             @                          �k@�E��ӭ�?             B@������������������������       �                     "@                          �b@��}*_��?             ;@������������������������       �R���Q�?             4@������������������������       �                     @                           �?*�8�4�?�            �k@                           �?��S���?'             N@                           �?<ݚ)�?             B@������������������������       �������?             .@������������������������       �                     5@                           �?      �?             8@������������������������       �                     2@������������������������       �      �?             @                          �e@ rc����?a            `d@                          �e@�p=
�c�?_             d@������������������������       ����7�?[            @c@������������������������       ��q�q�?             @              	          (33@�q�q�?             @������������������������       �                     �?������������������������       �                      @       .                    �?�Oܨ��?�            Pr@        '                    �J@�q�q�?A            �\@!       $                    �?ȵHPS!�?             J@"       #                   0j@�E��ӭ�?             2@������������������������       �                     @������������������������       ��r����?             .@%       &                   �d@г�wY;�?             A@������������������������       �                     �?������������������������       �                    �@@(       +                    q@�g�y��?"             O@)       *                    @ҳ�wY;�?             A@������������������������       ��<ݚ�?             ;@������������������������       �؇���X�?             @,       -                   �u@����X�?             <@������������������������       ��LQ�1	�?             7@������������������������       �                     @/       6                    �?x疑��?z            `f@0       3                    �?���c�H�?#            �H@1       2                   �q@      �?             @@������������������������       �                     =@������������������������       ��q�q�?             @4       5                    �?j���� �?             1@������������������������       �                     "@������������������������       �      �?              @7       :                    @$�q-�?W            @`@8       9                   @[@�f�¦ζ?F            �Z@������������������������       ��	j*D�?	             *@������������������������       ���K2��?=            �W@;       <                    �?��<b���?             7@������������������������       �X�Cc�?             ,@������������������������       �                     "@�t�bh�h(h+K ��h-��R�(KK=KK��ha�B�       @q@     0u@      k@     @Z@     �A@      P@      "@      K@      @      G@       @      A@      @      (@      @       @              @      @      @      :@      $@      "@              1@      $@      1@      @              @     �f@     �D@      @@      <@      &@      9@      &@      @              5@      5@      @      2@              @      @     �b@      *@     �b@      &@     `b@      @       @      @      �?       @      �?                       @     �M@     @m@      C@      S@      @      G@      @      *@      @               @      *@      �?     �@@      �?                     �@@      @@      >@      (@      6@      @      5@      @      �?      4@       @      4@      @              @      5@     �c@      &@      C@      �?      ?@              =@      �?       @      $@      @      "@              �?      @      $@      ^@      @     �Y@      @      "@      �?     @W@      @      2@      @      "@              "@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ9M�hG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK5hyh(h+K ��h-��R�(KK5��h��B�                             �?r�a����?�           8�@                           @|���>�?�            0w@       
       	          ���@�$�����?�            `n@                           �L@��Q�Vz�?�            �l@              	          033�?�fp�IЮ?g             d@������������������������       � � ���?e            �c@������������������������       ��q�q�?             @       	                    �M@H�V�e��?*             Q@������������������������       �X�<ݚ�?	             2@������������������������       �H%u��?!             I@                           �?d}h���?	             ,@                          �b@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                      @                           �?     ��?L             `@                           �?���Hx�?+             R@������������������������       �                     F@              
             �?      �?             <@������������������������       ����N8�?             5@������������������������       �؇���X�?             @                           �?������?!             L@                          �`@�*/�8V�?            �G@������������������������       �                     @������������������������       �&^�)b�?            �E@              	          ����?�<ݚ�?             "@������������������������       �                      @������������������������       �                     @       *       	          ����?<�'܀w�?�            �n@       #                    �?bf@����?8            �S@                            `@@�0�!��?             A@������������������������       �                     2@!       "                   @a@      �?             0@������������������������       �؇���X�?             @������������������������       �                     "@$       '                    @�q�q�?"            �F@%       &                    �?���@��?            �B@������������������������       ��t����?             1@������������������������       ��z�G��?             4@(       )                    �?      �?              @������������������������       �                     �?������������������������       �                     @+       0                   0b@|T(W�j�?f            �d@,       /                   �j@ �|ك�?J            �^@-       .                    @ qP��B�?            �E@������������������������       �                     E@������������������������       �                     �?������������������������       �        2             T@1       2                    �G@X�Cc�?             E@������������������������       �                      @3       4                   �n@�G�z�?             D@������������������������       �      �?             4@������������������������       �R���Q�?             4@�t�b��      h�h(h+K ��h-��R�(KK5KK��ha�BP       �r@     �s@     �\@     p@      >@     �j@      3@     @j@      @     �c@      @     `c@       @      �?      ,@      K@       @      $@      @      F@      &@      @      @      @              @      @               @              U@      F@     @P@      @      F@              5@      @      4@      �?      �?      @      3@     �B@      (@     �A@      @               @     �A@      @       @               @      @              g@     �M@      B@     �E@      @      <@              2@      @      $@      @      �?              "@      >@      .@      =@       @      .@       @      ,@      @      �?      @      �?                      @     �b@      0@     �^@      �?      E@      �?      E@                      �?      T@              ;@      .@               @      ;@      *@      $@      $@      1@      @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJpVhG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK3hyh(h+K ��h-��R�(KK3��h��B(                            Pb@ �����?�           8�@                           �?��M���?�            s@                           �?�S���,�?/            @T@              	          ���@`Ql�R�?            �G@������������������������       �                     G@������������������������       �                     �?       
                   �^@г�wY;�?             A@       	                   �]@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     >@                           @N@؇���X�?�             l@                          �e@�
�@c�?Z            �b@                          @Z@���;QU�?X            @b@������������������������       �                     �?������������������������       ���Ή�ν?W             b@������������������������       �                     @              	          ����?��{�?6�?.            �R@                           �?������?
             .@������������������������       �      �?              @������������������������       �                     @                          �`@�r����?$             N@������������������������       �                    �C@������������������������       ��ՙ/�?             5@       &       
             �?�C�^�?�            `s@       !                    �?��S���?C            @Z@                           @�L��7Q�?9            @V@                           �?j�q����?!             I@������������������������       ����Q��?             $@������������������������       �      �?             D@                            �O@��Sݭg�?            �C@������������������������       �b�h�d.�?            �A@������������������������       �                     @"       %                   pe@     ��?
             0@#       $                     @�8��8��?             (@������������������������       �                     �?������������������������       �                     &@������������������������       �                     @'       .                    �?�u�:T��?�            �i@(       +                    �?���+�?.            �R@)       *                    �?�G�5��?*            @Q@������������������������       �r�q��?%             N@������������������������       ��<ݚ�?             "@,       -       	          pff�?z�G�z�?             @������������������������       �                     @������������������������       �                     �?/       0                    @G@ �	.��?X            ``@������������������������       �                      H@1       2                   �b@�1/z��?8            �T@������������������������       �^l��[B�?*             M@������������������������       �                     9@�t�bh�h(h+K ��h-��R�(KK3KK��ha�B0       Ps@      s@     @l@     �S@      A@     �G@      �?      G@              G@      �?             �@@      �?      @      �?      @                      �?      >@              h@      @@      a@      *@      a@      $@              �?      a@      "@              @      L@      3@      @      &@      @      @              @      J@       @     �C@              *@       @     �T@     `l@     �H@      L@      C@     �I@      "@     �D@      @      @      @     �A@      =@      $@      =@      @              @      &@      @      &@      �?              �?      &@                      @      A@     `e@      5@     �J@      1@      J@      $@      I@      @       @      @      �?      @                      �?      *@     �]@              H@      *@     �Q@      *@     �F@              9@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ��hG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK/hyh(h+K ��h-��R�(KK/��h��BH
                             �?��>�'��?�           8�@              	          pff�?�&��?�             s@                           �?TV����?F            �]@                           @�p����?&            �N@                           �J@�[�IJ�?            �G@������������������������       �H%u��?             9@������������������������       ��GN�z�?             6@������������������������       �        	             ,@	                           �?�����?             �L@
                           b@�T|n�q�?            �E@������������������������       �ףp=
�?             D@������������������������       �                     @              	          ����?d}h���?	             ,@������������������������       �r�q��?             (@������������������������       �      �?              @                           @�*/�8V�?{            �g@              	          033�?����>�?/            �R@                           �?l��[B��?             =@������������������������       �ףp=
�?             $@������������������������       ��d�����?             3@                          �]@�����H�?            �F@������������������������       �        	             0@������������������������       �д>��C�?             =@������������������������       �        L            �\@       &                   �a@����2�?�            Ps@                          �j@B�
k���?'            �P@                           @�c�Α�?             =@                          Pc@���}<S�?             7@������������������������       �                      @������������������������       �                     5@������������������������       �                     @        #                    �?p�ݯ��?             C@!       "                    �?�eP*L��?             6@������������������������       �                      @������������������������       �؇���X�?	             ,@$       %                     R@      �?             0@������������������������       �؇���X�?             ,@������������������������       �                      @'       .                   `f@@1�`�?�            @n@(       +                    @�t����?�            �m@)       *                    �?���2"��?z             h@������������������������       �p��@���?j            @e@������������������������       ���<b���?             7@,       -                     D@��Hg���?#            �F@������������������������       �                      @������������������������       �RB)��.�?!            �E@������������������������       �                     @�t�bh�h(h+K ��h-��R�(KK/KK��ha�B�       �q@     �t@     �k@     �U@      J@     �P@      A@      ;@      4@      ;@      @      6@      1@      @      ,@              2@     �C@      @      B@      @      B@      @              &@      @      $@       @      �?      �?      e@      4@      K@      4@      ,@      .@      "@      �?      @      ,@      D@      @      0@              8@      @     �\@              P@     �n@      @@     �A@       @      5@       @      5@       @                      5@      @              8@      ,@      (@      $@               @      (@       @      (@      @      (@       @               @      @@     @j@      <@     @j@      1@      f@      (@     �c@      @      2@      &@      A@       @              "@      A@      @        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ��nhG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK!hyh(h+K ��h-��R�(KK!��h��B8                	          ����?Z�����?�           8�@                           �?�^���l�?9           @       
                   0f@�v:���?            �i@              	          pff�?     8�?u             h@                          @[@���0��?@             [@������������������������       �@�0�!��?             1@������������������������       �և���X�?8            �V@       	                   Pd@���H��?5             U@������������������������       �z�G�z�?             @������������������������       �l{��b��?2            �S@������������������������       �        
             (@                           @�2ن��?�            Pr@                           c@,��J�H�?�            @k@������������������������       �                      @                           �K@�`5���?�             k@������������������������       � g�yB�?X             `@������������������������       ������?8            �U@                           f@L�qA��?(            �R@              	             �?�iޤ��?$            �P@������������������������       ��b��[��?            �K@������������������������       ��8��8��?             (@������������������������       �                      @                           @�U�:��?P            �]@                           @�1�`jg�?J            �[@              	          `ff @�MI8d�?            �B@������������������������       �                      @                           �?(N:!���?            �A@������������������������       ����Q��?             $@������������������������       �                     9@������������������������       �        1            @R@               
             �?      �?              @������������������������       �                     @������������������������       �                     @�t�bh�h(h+K ��h-��R�(KK!KK��ha�B       �q@     �t@     @f@     �s@      `@     �R@      `@     �O@     �K@     �J@      @      ,@      J@     �C@     �R@      $@      �?      @     @R@      @              (@     �H@     �n@      5@     �h@       @              3@     �h@       @     �_@      1@     �Q@      <@     �G@      4@     �G@      3@      B@      �?      &@       @              [@      $@      Z@      @      ?@      @               @      ?@      @      @      @      9@             @R@              @      @              @      @        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJXk�hG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK)hyh(h+K ��h-��R�(KK)��h��B�                             �?��O���?�           8�@              	          pff�?�t����?�            �s@       
       	          833�?�r�����?L            @^@                          �c@�q�q�?2            �R@                          `c@6YE�t�?            �@@������������������������       ��GN�z�?             6@������������������������       �                     &@       	                    �?�G��l��?             E@������������������������       ��GN�z�?             6@������������������������       �R���Q�?             4@                          �m@�I� �?             G@������������������������       �        
             3@              
             �?X�<ݚ�?             ;@������������������������       �����X�?             5@������������������������       �                     @                           �Q@�C��2(�?~            �h@                          Pe@�}�+r��?z            �g@                          `a@@i�)ԙ�?s            �f@������������������������       � T���v�?E            @\@������������������������       �        .            @Q@                           @      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                      @                            @z�c�@-�?�            �r@                           c@�����?�            @j@������������������������       �                     @                           �K@ƺ"+L�?�            �i@������������������������       �        R            �`@                          �d@<ݚ�?2             R@������������������������       �Dc}h��?'             L@������������������������       �                     0@!       "                   @[@v ��?8            �U@������������������������       �                      @#       &                    �?�e����?3            �S@$       %                    _@     ��?             0@������������������������       �                     $@������������������������       �      �?             @'       (       
             �?�^�����?(             O@������������������������       �"Ae���?            �G@������������������������       ��r����?             .@�t�bh�h(h+K ��h-��R�(KK)KK��ha�B�       ps@      s@     �n@     �R@     @P@      L@      I@      9@      <@      @      1@      @      &@              6@      4@      @      1@      1@      @      .@      ?@              3@      .@      (@      .@      @              @     �f@      2@     �f@      $@     `f@      @     �[@      @     @Q@              �?      @              @      �?                       @     �P@     �l@      4@     �g@      @              1@     �g@             �`@      1@     �K@      1@     �C@              0@      G@      D@               @      G@      @@      *@      @      $@              @      @     �@@      =@      ?@      0@       @      *@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ0��JhG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK+hyh(h+K ��h-��R�(KK+��h��Bh	                             @:��au��?�           8�@              	          `ff @�4I�PJ�?�            Pw@                          `\@���Q��?�             t@������������������������       �                     1@                          �l@v�Mǔ�?�            �r@                           �?     p�?S             `@������������������������       �>A�F<�?             C@������������������������       �(;L]n�?:            �V@	       
                    �?>;�n�n�?u            �e@������������������������       �X�@��l�?]            �`@������������������������       ���]�T��?            �D@                          �e@f1r��g�?            �J@              
             �?�t����?            �I@                          �l@ףp=
�?             I@������������������������       ����N8�?             5@������������������������       �                     =@������������������������       �                     �?������������������������       �                      @       "                    �?�GN�z�?�            @n@                           �?8�$�>�?S             `@                           �?�q�q�?%             N@                          @[@     ��?             @@������������������������       �                     @������������������������       �X�Cc�?             <@                           @      �?             <@������������������������       �      �?
             0@������������������������       �      �?             (@                           �?�~t��?.            @Q@                           �?�7��?            �C@������������������������       �                     <@������������������������       �"pc�
�?             &@        !                    �L@������?             >@������������������������       �        	             .@������������������������       ���S���?
             .@#       $                   �Z@�=|+g��?K            @\@������������������������       �                     @%       (       
             �?�o�s(��?H            �[@&       '       	            �? }�Я��?8            @V@������������������������       �      �?             @������������������������       �        5            @U@)       *                     M@����X�?             5@������������������������       ���
ц��?
             *@������������������������       �                      @�t�bh�h(h+K ��h-��R�(KK+KK��ha�B�       `s@     s@     �^@     @o@     �S@     @n@      1@             �N@     @n@      $@     �]@      @      ?@      @     �U@     �I@      _@      9@     @[@      :@      .@     �F@       @     �F@      @     �F@      @      0@      @      =@                      �?               @     `g@     �K@      U@     �F@      9@     �A@      2@      ,@              @      2@      $@      @      5@      �?      .@      @      @     �M@      $@     �B@       @      <@              "@       @      6@       @      .@              @       @     �Y@      $@              @     �Y@      @      V@      �?      @      �?     @U@              .@      @      @      @       @        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJڡWhG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK5hyh(h+K ��h-��R�(KK5��h��B�                              �?����v��?�           8�@              	          033�?S:#��?�             v@       
                    �?��t��?�            �l@                           �?X�EQ]N�?�            �j@                           �?�~�4_��?6             V@������������������������       ������?             C@������������������������       ��:pΈ��?!             I@       	                   �^@,(��?L            �_@������������������������       �        $             N@������������������������       ��qM�R��?(            �P@              	          ����?��S���?             .@                           `@���Q��?             $@������������������������       �                     @������������������������       �                     @                           �I@z�G�z�?             @������������������������       �                     @������������������������       �      �?              @                           �?.T�߸��?M             _@                           �?����X�?4            @S@                           �?��
P��?            �A@������������������������       �        	             &@������������������������       ��q�q�?             8@                           �?�����?             E@������������������������       �؇���X�?             <@������������������������       �                     ,@                          �_@�*/�8V�?            �G@                           @X�Cc�?             ,@������������������������       �                     @������������������������       �                     "@                          �b@�C��2(�?            �@@������������������������       �z�G�z�?             .@������������������������       �        
             2@!       (                    �?(�`�F��?�            Pp@"       '       	          ����?x��-�?f            �c@#       &                   �c@�<ݚ�?            �F@$       %                    �K@�n_Y�K�?             :@������������������������       ��C��2(�?             &@������������������������       ����Q��?	             .@������������������������       �                     3@������������������������       �        J            �\@)       .       
             �?�7i���?B            �Y@*       +                    �?z�G�z�?             D@������������������������       �                     �?,       -       
             �?8�Z$���?            �C@������������������������       �                     @������������������������       ��8��8��?             B@/       2                    c@��a�n`�?(             O@0       1                    @4��?�?#             J@������������������������       ���<D�m�?             �H@������������������������       ��q�q�?             @3       4                    �?ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@�t�bh�h(h+K ��h-��R�(KK5KK��ha�BP       pr@      t@     �X@     �o@      @@     �h@      9@     �g@      3@     @Q@      (@      :@      @     �E@      @     @^@              N@      @     �N@      @       @      @      @      @                      @      �?      @              @      �?      �?     �P@     �L@     �K@      6@      1@      2@              &@      1@      @      C@      @      8@      @      ,@              (@     �A@      "@      @              @      "@              @      >@      @      (@              2@     �h@     @P@     �b@      $@     �A@      $@      0@      $@      $@      �?      @      "@      3@             �\@             �G@     �K@     �@@      @              �?     �@@      @              @     �@@      @      ,@      H@      @     �G@      @      G@       @      �?      "@      �?              �?      "@        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ:d�hG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK+hyh(h+K ��h-��R�(KK+��h��Bh	                             �?��S���?�           8�@                          Pb@J�4C��?�            �r@              	          pff�?@�qmNh�?k            `f@                           @I@�xGZ���?            �A@������������������������       �                     @                           �?J�8���?             =@������������������������       �                     @������������������������       ��q�q�?             8@	       
                    �?������?V             b@������������������������       �        5            �U@                           �Q@ 	��p�?!             M@������������������������       �h�����?             L@������������������������       �                      @                          0f@��0u���?N             ^@                          �d@*��ZE�?E            �Z@                           @�6����?2            @R@������������������������       �x�����?            �C@������������������������       �������?             A@                           �?"pc�
�?            �@@������������������������       �                     2@������������������������       ����Q��?             .@������������������������       �        	             ,@                            �?�� ��b�?�            �s@                           �?8�ƨxt�?�            �k@������������������������       �        5            @X@                          �p@���b��?Y             _@                           @ףp=
�?K             Y@������������������������       ��IєX�?5             Q@������������������������       �     ��?             @@                           �K@�q�q�?             8@������������������������       �                     @������������������������       �                     1@!       &                   �b@D�n�3�?;            �W@"       %       	          `ff�?�n_Y�K�?            �C@#       $       	          033�?���>4��?             <@������������������������       �8�A�0��?             6@������������������������       �                     @������������������������       �                     &@'       *                    �?����X�?#             L@(       )                   0d@П[;U��?             =@������������������������       �8�Z$���?             *@������������������������       �      �?
             0@������������������������       �                     ;@�t�bh�h(h+K ��h-��R�(KK+KK��ha�B�       �q@     �t@     �k@     �S@     �c@      4@      3@      0@              @      3@      $@              @      3@      @     �a@      @     �U@              K@      @      K@       @               @     �N@     �M@     �N@     �F@      A@     �C@       @      ?@      :@       @      ;@      @      2@              "@      @              ,@     �P@      o@      ;@     @h@             @X@      ;@     @X@      $@     �V@      @      P@      @      :@      1@      @              @      1@              D@     �K@      8@      .@      *@      .@      *@      "@              @      &@              0@      D@      0@      *@       @      &@      ,@       @              ;@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ�I]fhG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK+hyh(h+K ��h-��R�(KK+��h��Bh	                             �?��}��?x           8�@              	          033�?6�iL�?�             v@       
                    �?��x_F-�?�             s@                           �P@����X��?�            �n@                           @L@@݈g>h�?�            �l@������������������������       ��q�Y��?g            @e@������������������������       �д>��C�?!             M@       	                   �i@b�2�tk�?
             2@������������������������       �                     "@������������������������       ��<ݚ�?             "@              	          pff�?��S���?&             N@                          @i@�θ�?             :@������������������������       �                     @������������������������       ��C��2(�?             6@                          �\@������?             A@������������������������       �                     @������������������������       ��חF�P�?             ?@                           @M@      �?"             H@                           @�t����?             A@                           �?����X�?	             ,@������������������������       �                     @������������������������       ����Q��?             $@������������������������       �                     4@                          �h@և���X�?             ,@������������������������       �                     @                           �?�����H�?             "@������������������������       �                     @������������������������       ��q�q�?             @       $                    �?X�p���?�            Pp@       #                    @@i��M��?$            @P@                           �\@�iʫ{�?            �J@������������������������       �                     @!       "       	          033@H%u��?             I@������������������������       �=QcG��?            �G@������������������������       �                     @������������������������       �                     (@%       &                    �E@�[$�G�?z            �h@������������������������       �                      @'       (                   `@r ��*�?u            �g@������������������������       �                     @)       *       	          ����?�E��1�?s            �f@������������������������       �����X�?(            �O@������������������������       ��S���?K             ^@�t�bh�h(h+K ��h-��R�(KK+KK��ha�B�       0q@     @u@      X@      p@      N@     �n@      <@     @k@      5@     �i@      &@     �c@      $@      H@      @      &@              "@      @       @      @@      <@      @      4@      @               @      4@      :@       @              @      :@      @      B@      (@      >@      @      $@      @      @              @      @      4@              @       @      @              �?       @              @      �?       @     `f@     �T@      5@      F@      "@      F@      @              @      F@      @      F@      @              (@             �c@      C@               @     �c@      >@              @     �c@      9@     �F@      2@     @\@      @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ�޵#hG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK/hyh(h+K ��h-��R�(KK/��h��BH
                             �? �����?|           8�@                           �?�Pk���?�             y@       
                    @d/�@7�?S             a@                          �s@HP�s��?L            @_@                           @���U�?E            �\@������������������������       ��h����?D             \@������������������������       �                      @       	       	          ����?�eP*L��?             &@������������������������       �                     @������������������������       �                     @                           b@�q�q�?             (@������������������������       �                     @������������������������       �                      @              
             �?"X�8�?�            pp@              	          ����?��R[s�?G            @Z@                           @¦	^_�?             ?@������������������������       �                     (@������������������������       ��\��N��?             3@              
             �?,N�_� �?,            �R@������������������������       ��8��8��?             (@������������������������       �`Jj��?&             O@                           @L@"��S�&�?`            �c@                           @�S#א��?E            @]@������������������������       �@4և���?6            �X@������������������������       �p�ݯ��?             3@                          @k@D^��#��?            �D@������������������������       �@4և���?	             ,@������������������������       ��q�q�?             ;@       (                    �?6����?�            �j@       #                    �? 	��p�?l            �e@                           �Z@r�q��?)            �P@������������������������       �                      @!       "       	          ����?     ��?(             P@������������������������       �8�A�0��?             6@������������������������       �                     E@$       '                   �Z@`�߻�ɒ?C             [@%       &                    �?      �?             0@������������������������       �                     @������������������������       ��C��2(�?             &@������������������������       �        8             W@)       *                   �l@��]�T��?            �D@������������������������       �        
             4@+       .       
             �?����X�?             5@,       -                   �a@r�q��?
             2@������������������������       �                     &@������������������������       �և���X�?             @������������������������       �                     @�t�bh�h(h+K ��h-��R�(KK/KK��ha�B�        s@     Ps@      `@     �p@      2@     �]@      $@     �\@      @     �[@       @     �[@       @              @      @      @                      @       @      @              @       @             �[@      c@     �S@      ;@      "@      6@              (@      "@      $@     @Q@      @      &@      �?      M@      @     �@@     @_@      ,@     �Y@      @     �V@      @      (@      3@      6@      �?      *@      2@      "@      f@      C@     @d@      (@     �K@      &@               @     �K@      "@      *@      "@      E@             �Z@      �?      .@      �?      @              $@      �?      W@              .@      :@              4@      .@      @      .@      @      &@              @      @              @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ�G�hG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK)hyh(h+K ��h-��R�(KK)��h��B�                             @����v��?�           8�@              	          033�?��" ED�?�            �w@                           �?�]F���?�            t@                          �T@4�O)��?�            �n@������������������������       �                      @                           c@dLhg�?�            �n@������������������������       �0�N�]��?�            `l@������������������������       �b�2�tk�?	             2@	                           @P@      �?+            �R@
                           �?      �?              L@������������������������       ��C��2(�?            �@@������������������������       ���<b���?             7@                          Xq@�����H�?             2@������������������������       ��q�q�?             @������������������������       �                     (@                           @P̏����?%            �L@              
             �?@�0�!��?             �I@                          Ps@؇���X�?            �H@������������������������       �tk~X��?             B@������������������������       �                     *@������������������������       �                      @                           @O@r�q��?             @������������������������       �                     �?������������������������       �                     @       "       	          033�?l������?�            �m@              
             �?���>4��?4             U@������������������������       �                     @                          0m@X�<ݚ�?3            @T@                          �b@�������?             A@������������������������       �                     "@������������������������       ���H�}�?             9@        !                    [@��|�5��?            �G@������������������������       �                     @������������������������       �؇���X�?             E@#       (                   h~@�:�]��?`             c@$       '                    �?�.(�i��?_            �b@%       &                   �a@z�G�z�?&             I@������������������������       �                     4@������������������������       ��q�q�?             >@������������������������       �        9            @Y@������������������������       �                      @�t�bh�h(h+K ��h-��R�(KK)KK��ha�B�       pr@      t@     @[@     �p@     �P@     �o@      =@     @k@       @              ;@     @k@      4@     �i@      @      &@     �B@     �B@      5@     �A@      @      >@      2@      @      0@       @      @       @      (@             �E@      ,@      E@      "@      E@      @      =@      @      *@                       @      �?      @      �?                      @     @g@     �I@     �F@     �C@              @     �F@      B@      "@      9@              "@      "@      0@      B@      &@              @      B@      @     �a@      (@     �a@      $@      D@      $@      4@              4@      $@     @Y@                       @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ���JhG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK1hyh(h+K ��h-��R�(KK1��h��B�
                            �a@�.�t���?q           8�@       	                    �?�t�~U�?w            �f@                           �?b�2�tk�?             B@                           @>���Rp�?             =@                           �?��S���?
             .@������������������������       �      �?	             ,@������������������������       �                     �?������������������������       �                     ,@������������������������       �                     @
              	            �? )�y���?_             b@                          @j@     ��?             0@������������������������       �                     @                          �\@      �?	             (@������������������������       �                      @������������������������       �ףp=
�?             $@                           _@�7�	|��?S             `@������������������������       �        *            �O@                           @����e��?)            �P@������������������������       �$�q-�?	             *@������������������������       �                     �J@       $                    �?
�~z���?�             {@                           �?������?w            �h@                           �L@t�n_Y��?@             Z@                           @��.��?$            �N@������������������������       �                    �E@������������������������       �X�<ݚ�?             2@                          q@�+��<��?            �E@������������������������       ������?             5@������������������������       ��GN�z�?             6@       !                    @K@H~��D
�?7            �W@                            �H@8�A�0��?             6@������������������������       �                     @������������������������       �     ��?
             0@"       #                   �c@L������?)            @R@������������������������       ���s����?             E@������������������������       �                     ?@%       ,                    �?��k=.��?�            `m@&       )                    @�˹�m�?P             c@'       (                    �?@;�"�?A            �^@������������������������       �h�����?;             \@������������������������       ����|���?             &@*       +       
             �?8^s]e�?             =@������������������������       ���
ц��?             *@������������������������       �      �?	             0@-       .                    �H@j����?3            �T@������������������������       �                     1@/       0                    �?4���C�?(            �P@������������������������       ��q�q�?             B@������������������������       ��r����?             >@�t�bh�h(h+K ��h-��R�(KK1KK��ha�B       0s@     @s@     �c@      6@      6@      ,@      6@      @       @      @      @      @      �?              ,@                      @      a@       @      "@      @              @      "@      @               @      "@      �?      `@      �?     �O@             @P@      �?      (@      �?     �J@             �b@     �q@     �Y@      X@      =@     �R@      $@     �I@             �E@      $@       @      3@      8@       @      3@      1@      @     �R@      5@      "@      *@      @              @      *@     @P@       @      A@       @      ?@             �F@     �g@      1@     �`@       @     �\@      @      [@      @      @      "@      4@      @      @       @      ,@      <@     �K@              1@      <@      C@      8@      (@      @      :@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ�
HyhG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK7hyh(h+K ��h-��R�(KK7��h��B                
             �?��FY��?�           8�@                           @K@���-|$�?�            @s@              	          pff�?l��TO��?N            @_@                           �?�M;q��?.            �R@������������������������       �                     :@                           �?Tt�ó��?            �H@������������������������       ��	j*D�?             :@������������������������       ��㙢�c�?             7@	       
                   �i@H%u��?              I@������������������������       �                     4@                          �a@z�G�z�?             >@������������������������       �                     5@������������������������       ��q�q�?             "@                           �?2��7z��?x            �f@                           q@�f7�z�?(             M@                           �?�Gi����?            �B@������������������������       �                     @������������������������       �      �?             >@                           �N@�����?             5@������������������������       �        
             1@������������������������       �      �?             @                           �?h�N?���?P            @_@                           @ ��N8�?4             U@������������������������       �        3            �T@������������������������       �                     �?                           @���?            �D@������������������������       �     ��?             @@������������������������       ��<ݚ�?             "@       *                    @j�!����?�            0s@       %                   r@&!��Ji�?�            �n@       "       	          833�?     ��?x             h@        !       	          ����?�ص�ݒ�?R            @_@������������������������       �|�9ǣ�?M            �]@������������������������       �����X�?             @#       $                    �?0�,���?&            �P@������������������������       �                     �?������������������������       �����e��?%            �P@&       )                   u@H(���o�?             �J@'       (                   0e@��+��?            �B@������������������������       �d��0u��?             >@������������������������       �                     @������������������������       �        	             0@+       2                   �^@���@M^�?)             O@,       /                    �?�z�G��?             4@-       .                    Y@�t����?             1@������������������������       �                     @������������������������       �        	             (@0       1                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?3       4                    `@���N8�?             E@������������������������       �        	             1@5       6                    �?���Q��?             9@������������������������       ����y4F�?             3@������������������������       �                     @�t�bh�h(h+K ��h-��R�(KK7KK��ha�Bp       r@     `t@     �j@     �W@     �P@     �M@      6@     �J@              :@      6@      ;@      2@       @      @      3@      F@      @      4@              8@      @      5@              @      @     �b@     �A@      A@      8@      .@      6@              @      .@      .@      3@       @      1@               @       @     �\@      &@     �T@      �?     �T@                      �?      ?@      $@      =@      @       @      @     �R@      m@     �B@      j@      2@     �e@      0@     @[@      &@     �Z@      @       @       @     @P@      �?              �?     @P@      3@      A@      3@      2@      3@      &@              @              0@      C@      8@      @      ,@      @      (@      @                      (@      �?       @               @      �?              @@      $@      1@              .@      $@      .@      @              @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ���]hG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK1hyh(h+K ��h-��R�(KK1��h��B�
                             �?��a��?�           8�@              	          pff�?lD��+�?�            t@                           �?�ȋ}��?P            @`@              	            �?�2����?            �K@                          `i@�I�w�"�?             C@������������������������       �                     @������������������������       ���hJ,�?             A@������������������������       �                     1@	                           �?��H�}�?3            �R@
                           ]@d}h���?             E@������������������������       �        	             1@������������������������       ���H�}�?             9@                          0m@�eP*L��?            �@@������������������������       �      �?             4@������������������������       ��θ�?             *@                           @�g$����?q            �g@                           ^@:-�.A�?)            �P@������������������������       �                     :@              	          `ff
@D^��#��?            �D@������������������������       �d��0u��?             >@������������������������       �                     &@������������������������       �        H             _@       &                    @8RD�
��?�            `r@                          pc@<�����?�             i@                           �?�z�G��?5            �Q@                          �a@&y�X���?,             M@������������������������       �`2U0*��?             9@������������������������       �:ɨ��?            �@@                          �b@r�q��?	             (@������������������������       �                     @������������������������       �����X�?             @        #                    �?�Ώ��?V            ``@!       "                   �e@�J�T�?*            �Q@������������������������       �        %            �N@������������������������       �z�G�z�?             $@$       %                   �d@�8��8��?,             N@������������������������       ��q�q�?
             (@������������������������       �        "             H@'       *                   �a@�g�y��?7            @W@(       )                   �`@ףp=
�?             4@������������������������       �                     2@������������������������       �                      @+       .       	          pff�?��T���?*            @R@,       -                   q@tk~X��?             B@������������������������       �     ��?             @@������������������������       �                     @/       0                     I@��%��?            �B@������������������������       �                     "@������������������������       ���>4և�?             <@�t�bh�h(h+K ��h-��R�(KK1KK��ha�B       �r@     �s@     �l@      W@     �L@     @R@      "@      G@      "@      =@      @              @      =@              1@      H@      ;@     �@@      "@      1@              0@      "@      .@      2@      @      .@      $@      @     �e@      3@      H@      3@      :@              6@      3@      &@      3@      &@              _@             @R@     �k@      <@     �e@      5@     �H@      &@     �G@      �?      8@      $@      7@      $@       @      @              @       @      @      _@       @     @Q@             �N@       @       @      @     �K@      @      @              H@     �F@      H@      2@       @      2@                       @      ;@      G@      @      =@      @      =@      @              4@      1@      "@              &@      1@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ�;hG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK1hyh(h+K ��h-��R�(KK1��h��B�
                             @K@����v��?�           8�@                          �a@���>�?�            �r@                           @��ga�=�?+            �P@                           �?���|���?             6@������������������������       �        	             *@                           @J@�����H�?             "@������������������������       ��q�q�?             @������������������������       �                     @	       
       	          ����?����?�?            �F@������������������������       �                     �?������������������������       �                     F@                          pc@j(���?�            �l@                           �?�Z4���?*            �P@                           �H@��P���?            �D@������������������������       �և���X�?             5@������������������������       �                     4@                           \@�n_Y�K�?             :@������������������������       �                     @������������������������       �z�G�z�?             4@                           �?,���i�?h            �d@                           @t�e�í�?R            �`@������������������������       �        D            �[@������������������������       �\X��t�?             7@                           �?�q�q�?             >@������������������������       ����Q��?             9@������������������������       �                     @       &                    �?֕��9�?�            �s@       !       	          ���@�o+��?            �g@                          @W@�Q34�?l            �c@������������������������       �                     @                            i@�xO��(�?i             c@������������������������       �                     :@������������������������       ������?Y            �_@"       #                   `b@��a�n`�?             ?@������������������������       �                     8@$       %                     P@և���X�?             @������������������������       �                     @������������������������       �                     @'       ,       	          pff�?�N̸��?M            �_@(       +                   Pd@��R[s�?            �A@)       *                    [@�r����?             >@������������������������       �                     �?������������������������       �ܷ��?��?             =@������������������������       �                     @-       0                    @�nkK�?9             W@.       /                    �?��s����?             5@������������������������       ��X�<ݺ?             2@������������������������       �                     @������������������������       �        +            �Q@�t�bh�h(h+K ��h-��R�(KK1KK��ha�B       pr@      t@     @X@      i@      J@      .@       @      ,@              *@       @      �?       @      �?      @              F@      �?              �?      F@             �F@     @g@      9@      E@      "@      @@      "@      (@              4@      0@      $@              @      0@      @      4@      b@      $@      _@             �[@      $@      *@      $@      4@      $@      .@              @     �h@     �]@      U@     �Z@      L@     �Y@      @              I@     �Y@              :@      I@     @S@      <@      @      8@              @      @      @                      @     �\@      *@      :@      "@      :@      @              �?      :@      @              @      V@      @      1@      @      1@      �?              @     �Q@        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ� �thG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK1hyh(h+K ��h-��R�(KK1��h��B�
                             �?��}��?�           8�@                           @	�c��?            y@       
       	          ��� @�.�.���?�            Pq@                           �?(h�1W�?�            @p@                           @L@��0{9�?>            �W@������������������������       ����U�?&            �L@������������������������       �4�B��?            �B@       	                    @`�?�?n            �d@������������������������       ��#��g1�?h            �c@������������������������       ��<ݚ�?             "@                           @O@j���� �?             1@              	             
@�θ�?             *@������������������������       �                     @������������������������       �      �?              @������������������������       �                     @                           �?�d����?M            �^@                           �?H%u��?             I@                           @K@�q�q�?             (@������������������������       �                     @������������������������       �                     @                           �?P�Lt�<�?             C@������������������������       �                     9@������������������������       �$�q-�?	             *@                           �?�d�����?/            @R@                          �a@��Sݭg�?            �C@������������������������       ��q�q�?             "@������������������������       ��r����?             >@                           �?�!���?             A@������������������������       �     ��?             @@������������������������       �                      @       *                    �?�B�9ֆ�?�            �j@        %       	          pff�?�y��`�?i            �e@!       $                   Pd@d��0u��?!             N@"       #                    �?t�6Z���?            �K@������������������������       ����Q��?             $@������������������������       ��:�^���?            �F@������������������������       �                     @&       )                    �?�h����?H             \@'       (                   @i@�nkK�?             G@������������������������       ������?             5@������������������������       �                     9@������������������������       �        )            �P@+       ,                    �?^����?            �E@������������������������       �                     @-       .                   �l@>A�F<�?             C@������������������������       �        
             1@/       0                    @�q�q�?             5@������������������������       �                     *@������������������������       �      �?              @�t�bh�h(h+K ��h-��R�(KK1KK��ha�B       0q@     @u@     �Z@     `r@      =@      o@      3@      n@      ,@      T@       @     �K@      (@      9@      @      d@      @     @c@       @      @      $@      @      $@      @      @              @      @              @     @S@      G@      F@      @      @      @      @                      @     �B@      �?      9@              (@      �?     �@@      D@      $@      =@      @      @      @      :@      7@      &@      7@      "@               @      e@      G@     �c@      .@     �G@      *@     �G@       @      @      @     �D@      @              @     �[@       @      F@       @      3@       @      9@             �P@              (@      ?@      @              @      ?@              1@      @      ,@              *@      @      �?�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ��1hG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK3hyh(h+K ��h-��R�(KK3��h��B(                
             �?�������?�           8�@                           @H�g����?�            u@                          pb@����[��?d            �d@                          `d@��!pc�?7             V@������������������������       �                     @                           �?�<p���?3            �T@������������������������       ���ɉ�?)            @P@������������������������       �j���� �?
             1@	                           �?l������?-            �S@
              
             �?�\��N��?             3@������������������������       �                     @������������������������       �      �?
             0@                          `a@�r����?!             N@������������������������       ����.�6�?             G@������������������������       �X�Cc�?
             ,@                          �a@@�0�!��?l            @e@                          Xp@��:�-�??            @Y@������������������������       �                     �J@                          �p@ �q�q�?             H@������������������������       �                      @������������������������       �                     G@                          @d@��x�5��?-            @Q@              	          pff�?Rg��J��?"            �H@������������������������       ��KM�]�?             3@������������������������       ��z�G��?             >@              	          ����?ףp=
�?             4@������������������������       �r�q��?             (@������������������������       �                      @       (                    @����o�?�            `q@       #                    @L@H%u��?�             i@                            c@���N8�?P            �_@������������������������       �                     �?!       "                    �?`2U0*��?O            @_@������������������������       �`�(c�??            �X@������������������������       ��>����?             ;@$       %                   Pj@���"͏�?2            �R@������������������������       �        	             (@&       '                    �?¦	^_�?)             O@������������������������       �(N:!���?            �A@������������������������       �|��?���?             ;@)       0                    �L@      �?0            �S@*       -                    n@�J��%�?            �H@+       ,                   g@      �?             @@������������������������       �      �?             @������������������������       � ��WV�?             :@.       /                    c@�t����?             1@������������������������       �                     @������������������������       ��q�q�?             (@1       2                    @O@V�a�� �?             =@������������������������       �                     7@������������������������       �                     @�t�bh�h(h+K ��h-��R�(KK3KK��ha�B0       Pr@      t@     �l@     �Z@     �V@     @S@     @R@      .@              @     @R@      "@     �O@       @      $@      @      1@      O@      "@      $@      @              @      $@       @      J@      @     �E@      @      "@     �a@      >@     �X@       @     �J@              G@       @               @      G@             �D@      <@      7@      :@       @      1@      5@      "@      2@       @      $@       @       @             �O@     �j@      8@      f@      @      ^@      �?              @      ^@      @     �W@       @      9@      2@      L@              (@      2@      F@      @      ?@      ,@      *@     �C@     �C@      0@     �@@      @      <@      @      @      �?      9@      (@      @      @              @      @      7@      @      7@                      @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ�JIhG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK1hyh(h+K ��h-��R�(KK1��h��B�
                	          033�?���Y��?�           8�@                           @      �?�            �u@                          `\@h�3A_'�?�            pp@������������������������       �                     (@                          �r@���w;�?�            `o@                           �?d�cZյ�?�            �j@������������������������       ��# ��?x            �g@������������������������       �\X��t�?             7@	       
                    �?p9W��S�?             C@������������������������       ���� ��?             ?@������������������������       �                     @                           �?�Je\���?6            @T@                          �^@z�G�z�?             D@                           �G@r�q��?             @������������������������       �                     �?������������������������       �                     @                           �N@l��\��?             A@������������������������       ��g�y��?             ?@������������������������       ��q�q�?             @                           �?��P���?            �D@                           �L@H�V�e��?             A@������������������������       ��q�q�?             2@������������������������       �      �?	             0@                          @i@����X�?             @������������������������       �                     �?������������������������       �r�q��?             @       $                    @��M�?�            �p@       #       
             �?և���X�?P            �`@                            �?4=�%�?<            �X@              	          ���@�2�o�U�?#            �K@������������������������       ��*/�8V�?            �G@������������������������       �      �?              @!       "                    �O@Du9iH��?            �E@������������������������       �                     >@������������������������       ��θ�?             *@������������������������       �                    �A@%       ,                    �?���}<S�?Y            @a@&       )                    �? s�n_Y�?!             J@'       (                    �?�n_Y�K�?	             *@������������������������       �                     @������������������������       ������H�?             "@*       +       	          ����?$�q-�?            �C@������������������������       �z�G�z�?             $@������������������������       �XB���?             =@-       .                   �e@��f�{��?8            �U@������������������������       �        5            �T@/       0                   �j@�q�q�?             @������������������������       �                     �?������������������������       �                      @�t�bh�h(h+K ��h-��R�(KK1KK��ha�B       �p@     �u@     �U@      p@     �F@     @k@      (@             �@@     @k@      6@     �g@      "@     �f@      *@      $@      &@      ;@      @      ;@      @             �D@      D@      @@       @      �?      @      �?                      @      ?@      @      >@      �?      �?       @      "@      @@      @      ;@      @      (@      �?      .@       @      @      �?              �?      @     �f@      V@     �L@      S@     �L@     �D@      1@      C@      (@     �A@      @      @      D@      @      >@              $@      @             �A@     �_@      (@     �D@      &@      @       @      @              �?       @      B@      @       @       @      <@      �?     @U@      �?     �T@               @      �?              �?       @        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ��NhG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK)hyh(h+K ��h-��R�(KK)��h��B�                             @ד�w��?�           8�@                           �?f���?�            0v@              	          033�?      �?S            �_@                           �?��̅��?=            �W@              	          833�?P�%f��?:            �V@������������������������       �d�
��?             F@������������������������       ���<b���?             G@������������������������       �                     @	              
             �?��� ��?             ?@
                           �O@ףp=
�?             >@������������������������       �`2U0*��?             9@������������������������       ����Q��?             @������������������������       �                     �?                           �K@��F!�?�            �l@                           c@(;L]n�?c            �b@������������������������       �                      @              	          ����?PL��V�?b            �b@������������������������       � 7���B�?:            @T@������������������������       �        (            �P@                           @N@�6i����?0            �S@                           �?�G�z��?             D@������������������������       �r�q��?             8@������������������������       �      �?             0@������������������������       �                    �C@                          @[@&����?�            @p@                          0m@�8��8��?             (@������������������������       �                     @                          �m@r�q��?             @������������������������       �                     �?������������������������       �                     @       $                    �?ڏ�&��?�             o@        #       	          ����?�1��?o            �e@!       "                   ``@tk~X��?             B@������������������������       ������?             5@������������������������       ��q�q�?             .@������������������������       �        X             a@%       &                   `\@�EH,���?2            �R@������������������������       �                     $@'       (       	          pff�?�G\�c�?-            @P@������������������������       �     ��?             0@������������������������       ��J��%�?!            �H@�t�b�6     h�h(h+K ��h-��R�(KK)KK��ha�B�        r@     Pt@     �U@     �p@     �O@     �O@      B@     �M@      ?@     �M@      5@      7@      $@      B@      @              ;@      @      ;@      @      8@      �?      @       @              �?      7@     �i@      @      b@       @              @      b@      @     �S@             �P@      2@     �N@      2@      6@      @      4@      ,@       @             �C@     �i@      L@      �?      &@              @      �?      @      �?                      @     `i@     �F@     �d@      @      =@      @      3@       @      $@      @      a@             �B@      C@      $@              ;@      C@      &@      @      0@     �@@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ2�3hG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK5hyh(h+K ��h-��R�(KK5��h��B�                             �?�p ��?}           8�@                           �?~��D�?�            py@       
       	          ���@R��O��?�            pp@                           �?��)���?�            `o@                          �`@`�(c�?             �H@������������������������       ��xGZ���?            �A@������������������������       �                     ,@       	                    @x�7Fb��?z            @i@������������������������       ���8=��?a            �d@������������������������       �p�ݯ��?             C@                           @�q�q�?             (@������������������������       �                     @                          �d@և���X�?             @������������������������       �                     @������������������������       �                     @                           @H@�q�q�?^             b@                           �?�X�<ݺ?             2@                           �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        
             0@                           �?���f��?R            �_@              	          ����?��مD�?2            @S@������������������������       �      �?             >@������������������������       �`�q�0ܴ?            �G@                           @O@Rg��J��?             �H@������������������������       �     ��?             @@������������������������       ��t����?             1@       &                    �I@0��k���?~             j@       %                   �n@�q�q�?             H@       "                    @F@f���M�?             ?@        !                    m@r�q��?	             (@������������������������       ��C��2(�?             &@������������������������       �                     �?#       $                    �?�}�+r��?             3@������������������������       �؇���X�?             @������������������������       �                     (@������������������������       �                     1@'       .                    �?\���(\�?_             d@(       +                    �?��U/��?"            �L@)       *                    @O@���N8�?             5@������������������������       �        
             0@������������������������       �z�G�z�?             @,       -                    �?X�<ݚ�?             B@������������������������       �      �?             0@������������������������       ��z�G��?
             4@/       2                    �O@X�?٥�?=            �Y@0       1                    �?����ȫ�?1            �T@������������������������       �        +            �Q@������������������������       ��C��2(�?             &@3       4                    �?��s����?             5@������������������������       �z�G�z�?             @������������������������       �                     0@�t�bh�h(h+K ��h-��R�(KK5KK��ha�BP       �r@     �s@     �`@     q@      I@     �j@      E@      j@      3@      >@      3@      0@              ,@      7@     `f@      "@     `c@      ,@      8@       @      @      @              @      @      @                      @      U@      N@      �?      1@      �?      �?      �?                      �?              0@     �T@     �E@      N@      1@      .@      .@     �F@       @      7@      :@      5@      &@       @      .@     �d@      E@      <@      4@      &@      4@      $@       @      $@      �?              �?      �?      2@      �?      @              (@      1@             @a@      6@      D@      1@      4@      �?      0@              @      �?      4@      0@      ,@       @      @      ,@     �X@      @     @T@      �?     �Q@              $@      �?      1@      @      �?      @      0@        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJk�ahG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK-hyh(h+K ��h-��R�(KK-��h��B�	                	          033�?���i��?�           8�@                           �?�ⶕ��?0           P}@       
                    @���Q��?            `h@                           �?f<t=9%�?B             [@                            N@�7�QJW�?-            �R@������������������������       �                      J@������������������������       �\X��t�?             7@       	       	          ����?6YE�t�?            �@@������������������������       �     ��?
             0@������������������������       �                     1@                           �O@�=C|F�?=            �U@                           �M@,N�_� �?5            �R@������������������������       �6uH���?+             O@������������������������       �        
             (@                          (p@��
ц��?             *@������������������������       ��<ݚ�?             "@������������������������       �                     @                          �d@��t�0�?�             q@                           @��C�iF�?j            �e@                          �l@&��f���?\            @b@������������������������       � 7���B�?              K@������������������������       �8����?<             W@                           o@|��?���?             ;@������������������������       �@4և���?             ,@������������������������       �                     *@                          �e@T��,��?G            @Y@                          �[@`�LVXz�?E            �X@������������������������       ������H�?             "@������������������������       �        A            �V@������������������������       �                      @       *       
             �?��ӄ���?^            @b@        '                   �e@$�q-�?R            @`@!       $       
             �?������?M            �^@"       #                   �k@\-��p�?             =@������������������������       �                     *@������������������������       �      �?             0@%       &                    �N@`Ql�R�?9            �W@������������������������       �        ,            �Q@������������������������       ����}<S�?             7@(       )                    @և���X�?             @������������������������       �                     @������������������������       �                     @+       ,                    @     ��?             0@������������������������       �                     "@������������������������       �                     @�t�bh�h(h+K ��h-��R�(KK-KK��ha�B�       0r@     @t@     �d@     s@     @]@     �S@     �D@     �P@      *@      O@              J@      *@      $@      <@      @      &@      @      1@              S@      &@     @Q@      @     �L@      @      (@              @      @      @       @              @     �G@     `l@      F@      `@      >@      ]@       @      J@      <@      P@      ,@      *@      �?      *@      *@              @     �X@      �?     �X@      �?       @             �V@       @             �_@      3@      ^@      $@     @]@      @      9@      @      *@              (@      @      W@       @     �Q@              5@       @      @      @      @                      @      @      "@              "@      @        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ6ޤhG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK1hyh(h+K ��h-��R�(KK1��h��B�
                             �?BM�e�x�?           8�@                           @M@��Iߪ��?�            �w@                           �?ޅ��Rz�?�            �q@                           �?0?R����?�            �j@������������������������       �        -            @T@              	          033�?6YE�t�?V            �`@������������������������       ��C��2(�?P            @^@������������������������       �"pc�
�?             &@	                           �?&ջ�{��?%            @R@
                           @��h!��?            �L@������������������������       ���
ц��?             :@������������������������       �`Jj��?             ?@������������������������       �                     0@                          �p@�P�*�?8            @W@                          a@����X�?&            �Q@                          pb@p�ݯ��?
             3@������������������������       �      �?	             0@������������������������       �                     @                          0c@>a�����?            �I@������������������������       �r֛w���?             ?@������������������������       �        	             4@                          a@�㙢�c�?             7@                          ps@      �?             @������������������������       �                      @������������������������       �                      @                           @O@�KM�]�?             3@������������������������       �        
             .@������������������������       �      �?             @       "                    @F@�k��(A�?�            �m@       !                   �\@@4և���?             ,@                            �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     "@#       *       	          033�?��%����?�            �k@$       '                    �?
;&����?@             W@%       &                   �Z@����>�?            �B@������������������������       �                     @������������������������       �"pc�
�?            �@@(       )                    �?�2�o�U�?'            �K@������������������������       �                     @������������������������       ����c�H�?$            �H@+       .       	          ����?����?T            @`@,       -       
             �?�����H�?!             K@������������������������       ��nkK�?             G@������������������������       �      �?              @/       0       	          `ff @�"w����?3             S@������������������������       ��}�+r��?             3@������������������������       �        &            �L@�t�bh�h(h+K ��h-��R�(KK1KK��ha�B       �p@     �u@      Y@     pq@     �N@      l@      4@      h@             @T@      4@      \@      &@     �[@      "@       @     �D@      @@     �D@      0@      (@      ,@      =@       @              0@     �C@      K@      4@      I@      (@      @      (@      @              @       @     �E@       @      7@              4@      3@      @       @       @       @                       @      1@       @      .@               @       @      e@      Q@      �?      *@      �?      @      �?                      @              "@     �d@     �K@      F@      H@      ;@      $@              @      ;@      @      1@      C@      @              &@      C@     �^@      @      H@      @      F@       @      @      @     �R@      �?      2@      �?     �L@        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ��{hG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK-hyh(h+K ��h-��R�(KK-��h��B�	                            pb@*�3�V��?s           8�@                           �?��h!��?�            �q@              	          pff�?6�\"���?L            �_@                           �K@>a�����?            �I@������������������������       �                     B@              	          @33�?��S���?
             .@������������������������       ����Q��?             $@������������������������       �z�G�z�?             @	                           @�=A�F�?.             S@
                           �?      �?             :@������������������������       �     ��?	             0@������������������������       �                     $@                          �d@`2U0*��?             I@������������������������       �                     H@������������������������       �                      @              
             �?p#�����?`            �c@                           �?Tۢ��(�?P            �`@                           @���B���?              J@������������������������       �؇���X�?            �H@������������������������       �                     @                          �p@��'�`�?0            �T@������������������������       ��?�|�?            �B@������������������������       �                     G@                          �j@
;&����?             7@������������������������       �                     &@                           �?�8��8��?             (@������������������������       �                     @������������������������       �؇���X�?             @       ,       	          ���@�1�`jg�?�            �t@       %                    �?���@;��?�            �s@       "                    �?\�����?>            �[@        !                   Hq@���-T��?$             O@������������������������       �����?�?            �F@������������������������       ���.k���?             1@#       $                    �?8��8���?             H@������������������������       �д>��C�?             =@������������������������       �                     3@&       )       
             �?���`L�?�            �i@'       (                   �b@Z�K�D��?!            �G@������������������������       ����!pc�?             &@������������������������       �      �?             B@*       +                    @L@p=
ףp�?a             d@������������������������       ��h����?C             \@������������������������       �      �?             H@������������������������       �                     *@�t�bh�h(h+K ��h-��R�(KK-KK��ha�B�       �r@     �s@     �i@      T@     @Q@      M@       @     �E@              B@       @      @      @      @      @      �?     �N@      .@      *@      *@      *@      @              $@      H@       @      H@                       @      a@      6@      _@      &@      E@      $@      E@      @              @     �T@      �?      B@      �?      G@              (@      &@      &@              �?      &@              @      �?      @      X@     @m@     �T@     @m@      J@      M@      "@     �J@      �?      F@       @      "@     �E@      @      8@      @      3@              ?@      f@      1@      >@       @      @      "@      ;@      ,@     @b@       @     �[@      (@      B@      *@        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ?{�hG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK1hyh(h+K ��h-��R�(KK1��h��B�
                             @K@j�[.��?�           8�@              	          033�?���-|$�?�            @s@                           �?�|�
��?�            �o@������������������������       �        3            �T@              
             �?'��%��?k            �e@                           �?֭��F?�?            �G@������������������������       �$��m��?             :@������������������������       ����N8�?             5@	       
                    c@6C�d�?L            �_@������������������������       �                      @������������������������       � E=��H�?K             _@                           �?^�!~X�?!            �J@                            G@�q�q�?	             (@������������������������       �                     @������������������������       �                      @                           @F@��p\�?            �D@������������������������       �                     8@                          �`@@�0�!��?             1@������������������������       �                     $@������������������������       �և���X�?             @       $       	          `ff�?b��W��?�            0s@                           �?����p�?_             a@                           @R=6�z�?.            @P@                           �L@      �?&             L@������������������������       ���.k���?
             1@������������������������       ��ݜ�?            �C@                           �M@X�<ݚ�?             "@������������������������       �                     @������������������������       �                     @       !                    �?R_u^|�?1            �Q@                           `b@�eP*L��?              F@������������������������       �                      @������������������������       �X�<ݚ�?             B@"       #                    [@������?             ;@������������������������       �                     @������������������������       �                     4@%       *                    �?J��$���?k            `e@&       '                    ]@�e�,��?%            �M@������������������������       �                     @(       )                    �L@�c�����?             �J@������������������������       �      �?             ,@������������������������       �8�Z$���?            �C@+       .       
             �?      �?F             \@,       -                    �?`�E���?>            @X@������������������������       �        '            @Q@������������������������       �@4և���?             <@/       0                    `P@�q�q�?             .@������������������������       �                     $@������������������������       �                     @�t�bh�h(h+K ��h-��R�(KK1KK��ha�B       �r@     �s@     �W@     �j@      H@     �i@             �T@      H@     @_@      =@      2@      "@      1@      4@      �?      3@     �Z@       @              1@     �Z@      G@      @       @      @              @       @              C@      @      8@              ,@      @      $@              @      @     �i@     �Y@     �M@     @S@      3@      G@      ,@      E@      "@       @      @      A@      @      @      @                      @      D@      ?@      4@      8@               @      4@      0@      4@      @              @      4@              b@      :@      D@      3@              @      D@      *@      @      @     �@@      @     @Z@      @     �W@       @     @Q@              :@       @      $@      @      $@                      @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ��}whG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK;hyh(h+K ��h-��R�(KK;��h��B�                            Pb@ד�w��?y           8�@                           �O@Ɔdq��?�            `q@       
                    �?�8=�?~            �i@                          @\@�8��8��?Z             b@                           ^@      �?             8@������������������������       �                     "@������������������������       ����Q��?
             .@       	                    @�(\����?K             ^@������������������������       ��˹�m��?             C@������������������������       �        4            �T@                           _@`՟�G��?$             O@                          �X@؇���X�?             <@������������������������       �                      @������������������������       �$�q-�?             :@                           �?�t����?             A@������������������������       �"pc�
�?             6@������������������������       �      �?             (@              	          ����?�q�q�?%             R@                           �P@�>����?             ;@                           @z�G�z�?             $@������������������������       �                      @������������������������       �                      @������������������������       �                     1@                           ]@F�����?            �F@                          @Z@@4և���?             ,@������������������������       �                     �?������������������������       �                     *@                           �?��� ��?             ?@������������������������       ��q�q�?             @������������������������       �                     9@       ,                    �?��疾�?�            u@        '                    �?��B����?D             Z@!       $                    �? ��*��?>            �W@"       #       	          ����?��$�4��?%            �M@������������������������       �"pc�
�?"            �K@������������������������       �      �?             @%       &                    �L@�#-���?            �A@������������������������       �      �?
             (@������������������������       �                     7@(       )       
             �?ףp=
�?             $@������������������������       �                     @*       +                    \@�q�q�?             @������������������������       �                     �?������������������������       �                      @-       4                    @8ӈ(�3�?�             m@.       1                    @L@،c�u��?r             g@/       0                   @[@h�����?Y            �a@������������������������       ��n_Y�K�?             *@������������������������       �        R            �_@2       3                   @a@f.i��n�?            �F@������������������������       ��	j*D�?             *@������������������������       �     ��?             @@5       8       	          ����?     ��?              H@6       7                    �?@4և���?             ,@������������������������       �                     $@������������������������       �      �?             @9       :                    �?j���� �?             A@������������������������       ���X��?             <@������������������������       �r�q��?             @�t�bh�h(h+K ��h-��R�(KK;KK��ha�B�        r@     Pt@     �h@     �T@     �d@      D@     �`@      (@      .@      "@      "@              @      "@     @]@      @     �A@      @     �T@              A@      <@      8@      @               @      8@       @      $@      8@      @      2@      @      @      >@      E@       @      9@       @       @       @                       @              1@      <@      1@      �?      *@      �?                      *@      ;@      @       @      @      9@             �W@     `n@      K@      I@     �F@     �H@      *@      G@      $@     �F@      @      �?      @@      @      "@      @      7@              "@      �?      @               @      �?              �?       @              D@      h@      3@     �d@      @     �`@      @       @             �_@      ,@      ?@      "@      @      @      ;@      5@      ;@      �?      *@              $@      �?      @      4@      ,@      3@      "@      �?      @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ�,�hG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK3hyh(h+K ��h-��R�(KK3��h��B(                             �?T�h��?�           8�@                           �?���U��?�             s@                           �?      �?U             _@                          @e@     ��?-             P@                           �?�7����?"            �G@������������������������       ��C��2(�?             6@������������������������       �� �	��?             9@������������������������       �                     1@	                           [@���*�?(             N@
              	          ����?      �?              @������������������������       �                     @������������������������       �                     @                           �L@ȵHPS!�?#             J@������������������������       �      �?	             (@������������������������       ���(\���?             D@                           @<�Z��?g            �f@                          `b@�G�z.�?0             T@������������������������       �        $             L@                           �?�q�q�?             8@������������������������       �P���Q�?	             4@������������������������       �                     @              	          ����?`2U0*��?7             Y@                           �?�q�q�?
             (@������������������������       �؇���X�?             @������������������������       ����Q��?             @������������������������       �        -             V@       $                   �a@��\ck�?�            ps@       #       	          `ff�?��S���?$             N@                            �?���Q �?            �H@                          �^@��Q��?             4@������������������������       �                     @������������������������       �j���� �?	             1@!       "                   �o@\-��p�?             =@������������������������       �                     5@������������������������       �      �?              @������������������������       �                     &@%       ,                    �?@��:���?�            `o@&       )       
             �?4�0_���?�            @l@'       (                    �?b:�&���?5            �T@������������������������       �                     =@������������������������       ��E��ӭ�?#             K@*       +                    �?p�[&�?W            �a@������������������������       �                      H@������������������������       ��==Q�P�?7            �W@-       0                    a@�q�����?             9@.       /                    �?�θ�?
             *@������������������������       �                     @������������������������       ��z�G��?             $@1       2                    o@r�q��?
             (@������������������������       �                     "@������������������������       ��q�q�?             @�t�bh�h(h+K ��h-��R�(KK3KK��ha�B0       Pq@      u@     `k@     @U@      O@      O@      *@     �I@      *@      A@       @      4@      &@      ,@              1@     �H@      &@      @      @      @                      @      G@      @      "@      @     �B@      @     �c@      7@     �N@      3@      L@              @      3@      �?      3@      @              X@      @       @      @      @      �?       @      @      V@              M@     �o@      <@      @@      1@      @@      *@      @      @              $@      @      @      9@              5@      @      @      &@              >@     �k@      2@      j@      .@      Q@              =@      .@     �C@      @     �a@              H@      @      W@      (@      *@      $@      @      @              @      @       @      $@              "@       @      �?�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ�%\hG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK5hyh(h+K ��h-��R�(KK5��h��B�                             @���i��?w           8�@              	          033�?�l��� �?�            �x@                           �?Tpƥ��?�            `t@                           �?�IєX�?_             c@                          c@ףp=
�?8            �V@������������������������       �z�G�z�?             >@������������������������       �P���Q�?$             N@������������������������       �        '            �O@	                           �?��R�(��?b            �e@
                          0f@�G�z��?              N@������������������������       ����j��?             G@������������������������       �        
             ,@                           �?��(�?B            @\@������������������������       ��n_Y�K�?             *@������������������������       �HP�s��?:             Y@                           d@�㙢�c�?'            @Q@                           @O@X��Oԣ�?"             O@                          pb@�nkK�?             G@������������������������       �                     <@������������������������       ������H�?             2@                          Pn@     ��?	             0@������������������������       ��q�q�?             @������������������������       �ףp=
�?             $@              	          ����?����X�?             @������������������������       �                      @������������������������       �                     @       (                    �?ƯsY�h�?�            �k@       !                   �^@��.���?8            �U@               	          ����?���Q��?             9@                          �e@      �?
             0@������������������������       �                     �?������������������������       �        	             .@������������������������       �                     "@"       %                    d@ƆQ����?&            �N@#       $       	            �?8��8���?             H@������������������������       ����|���?             &@������������������������       ��?�|�?            �B@&       '                    �I@�	j*D�?             *@������������������������       ��q�q�?             @������������������������       �                     @)       0       	          833�?�qM�R��?W            �`@*       -                    @�θ�?            �C@+       ,                   @X@��hJ,�?             A@������������������������       �                     @������������������������       �`Jj��?             ?@.       /                   �`@z�G�z�?             @������������������������       �                     @������������������������       �                     �?1       4       	          ����?�==Q�P�?>            �W@2       3                    @��(\���?             D@������������������������       �Pa�	�?            �@@������������������������       �����X�?             @������������������������       �        #            �K@�t�bh�h(h+K ��h-��R�(KK5KK��ha�BP       0r@     @t@      \@     �q@     �K@     �p@      "@      b@      "@     @T@      @      8@      @     �L@             �O@      G@     �_@     �@@      ;@     �@@      *@              ,@      *@      Y@      @       @       @      W@     �L@      (@     �K@      @      F@       @      <@              0@       @      &@      @       @      @      "@      �?       @      @       @                      @     `f@     �D@     �L@      =@      $@      .@      �?      .@      �?                      .@      "@             �G@      ,@     �E@      @      @      @      B@      �?      @      "@      @       @              @     �^@      (@      >@      "@      =@      @              @      =@       @      �?      @              @      �?              W@      @     �B@      @      @@      �?      @       @     �K@        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ2�hG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK7hyh(h+K ��h-��R�(KK7��h��B                            Pb@r � 	��?�           8�@                           �?��O�;��?�             p@                           �?�6Re�?q            `f@                          �]@X�Emq�?$            �J@������������������������       �        
             .@                           @\�Uo��?             C@������������������������       �     ��?             @@������������������������       �                     @	                           �?�i�y�?M            �_@
                           �?��:x�ٳ?:            �X@������������������������       �        $            �P@������������������������       �      �?             @@������������������������       �                     ;@                           @���/��?4            �S@                           a@���|���?             F@              	          ����?��S���?             >@������������������������       �                     $@������������������������       ��z�G��?             4@                            N@؇���X�?             ,@������������������������       ��q�q�?             @������������������������       �                      @                           _@<=�,S��?            �A@������������������������       �                     .@              	          ����?��Q��?             4@������������������������       �                     @������������������������       �      �?	             ,@       (                    @���W!h�?�            Pv@       !                    �?|�(��?�            �o@                            �?     ��?>             X@                          `a@�+e�X�?2            �R@������������������������       ��2����?%            �K@������������������������       ��G�z��?             4@������������������������       �                     5@"       %                   �t@�7��?Y            �c@#       $                    �?��<�Ұ?T            `b@������������������������       ��Μ�5�?>            �[@������������������������       ��8��8��?             B@&       '                   d@�q�q�?             "@������������������������       �                     @������������������������       �                     @)       0                    �L@և���X�?H            @Z@*       -       
             �?�E��
��?'             J@+       ,                   �m@d}h���?             ,@������������������������       �                      @������������������������       �      �?             @.       /                    �?�d�����?             C@������������������������       �$�q-�?             :@������������������������       ��q�q�?             (@1       4                    @Ȩ�I��?!            �J@2       3                    �P@�㙢�c�?             G@������������������������       ��FVQ&�?            �@@������������������������       ���
ц��?             *@5       6                   �c@؇���X�?             @������������������������       �                     @������������������������       �                     �?�t�bh�h(h+K ��h-��R�(KK7KK��ha�Bp       @q@     0u@     �g@      Q@      c@      ;@      >@      7@      .@              .@      7@      "@      7@      @             �^@      @     �W@      @     �P@              <@      @      ;@              C@     �D@      0@      <@      ,@      0@              $@      ,@      @       @      (@       @      @               @      6@      *@      .@              @      *@              @      @      @     �U@     �p@      :@     @l@      2@     �S@      2@     �L@      "@      G@      "@      &@              5@       @     �b@      @     �a@       @     @[@      @     �@@      @      @      @                      @      N@     �F@      5@      ?@      &@      @       @              @      @      $@      <@       @      8@       @      @     �C@      ,@      C@       @      ?@       @      @      @      �?      @              @      �?        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ��(.hG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK/hyh(h+K ��h-��R�(KK/��h��BH
                            pb@ �����?�           8�@              
             �?f	���?�            0q@       
                    �?���^�?�            �k@                           @��ɹ?r            �g@                           �?�t����?,             Q@������������������������       ��(\����?             D@������������������������       �      �?             <@       	                    �? �.�?Ƞ?F             ^@������������������������       �        &            @P@������������������������       �h㱪��?             �K@                           �?�xGZ���?            �A@������������������������       �                     @              	            �?d��0u��?             >@������������������������       �                     @������������������������       �R�}e�.�?             :@                          �c@���3�E�?             J@                           �?�-���?             I@������������������������       �                     8@                          �n@      �?             :@������������������������       ���Q��?             4@������������������������       �                     @������������������������       �                      @       $                    �?@�ܻ��?�            @u@                          �d@؇���X�?�             l@                           �?�q-�?�             j@                           @���X�?$             L@������������������������       ���(\���?             D@������������������������       �      �?             0@                           \@`-�I�w�?b             c@������������������������       ��q�q�?             .@������������������������       ����Z�?W             a@        !                    �?     ��?
             0@������������������������       �                     @"       #       	          ����?��
ц��?             *@������������������������       ��q�q�?             "@������������������������       �                     @%       (                   �h@��o	��?L             ]@&       '                    �?@4և���?             ,@������������������������       �                     �?������������������������       �                     *@)       ,                    @$ޗQ��?D            �Y@*       +                   �\@�q�q�?$            �L@������������������������       �z�G�z�?             $@������������������������       ���|�5��?            �G@-       .                    �P@��S�ۿ?             �F@������������������������       � qP��B�?            �E@������������������������       �                      @�t�bh�h(h+K ��h-��R�(KK/KK��ha�B�        s@     Ps@     �j@     �O@     �h@      :@     @f@      $@      N@       @     �C@      �?      5@      @     �]@       @     @P@             �J@       @      3@      0@              @      3@      &@              @      3@      @      .@     �B@      *@     �B@              8@      *@      *@      @      *@      @               @             �W@     �n@      @@      h@      9@     �f@      .@     �D@      @     �B@      (@      @      $@     �a@      @      $@      @     �`@      @      "@              @      @      @      @      @      @              O@      K@      �?      *@      �?                      *@     �N@     �D@      3@      C@       @       @      &@      B@      E@      @      E@      �?               @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJx�+hG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK-hyh(h+K ��h-��R�(KK-��h��B�	                	          033�?�:�Ӛ��?�           8�@                           @(���@��?0           `}@       
                    �?F.< ?�?�            �t@                           �?ԼI�5��?�            �p@                           �?�C+����?C            @Y@������������������������       � ��~���??            �V@������������������������       �"pc�
�?             &@       	                   �m@�k2;���?m            �d@������������������������       �        >             V@������������������������       �p`q�q��?/            �S@                           �?�P�*�?%             O@                          �b@�5��
J�?             G@������������������������       �$G$n��?            �B@������������������������       ��q�q�?             "@              	          ����?      �?             0@������������������������       �r�q��?             @������������������������       �                     $@                           �O@��>4և�?[            �a@                           �?�������?N             ]@                          �m@8�Z$���?4            �S@������������������������       �^������?            �A@������������������������       �                     �E@                          �a@\�Uo��?             C@������������������������       �                     @������������������������       �:ɨ��?            �@@                          Pd@r�q��?             8@                          pk@�C��2(�?             6@������������������������       �      �?              @������������������������       �P���Q�?	             4@������������������������       �                      @                           �Z@ Ϸ�~�?X             b@������������������������       �                     �?!       &                   �a@�����H�?W             b@"       %                    @��F�D�?:            �X@#       $                    �? �#�Ѵ�?            �E@������������������������       ��q�q�?             @������������������������       ��(\����?             D@������������������������       �        "             L@'       *       	          033@f.i��n�?            �F@(       )                   @_@      �?             0@������������������������       �      �?              @������������������������       �      �?              @+       ,                   @n@\-��p�?             =@������������������������       �                     5@������������������������       �      �?              @�t�bh�h(h+K ��h-��R�(KK-KK��ha�B�       `q@     u@     �b@      t@     @P@     �p@      =@     �m@      6@     �S@      *@     @S@      "@       @      @      d@              V@      @      R@      B@      :@     �A@      &@      @@      @      @      @      �?      .@      �?      @              $@     @U@     �K@     @T@     �A@     �P@      (@      7@      (@     �E@              .@      7@      @              $@      7@      @      4@       @      4@      �?      �?      �?      3@       @              `@      1@              �?      `@      0@     @X@       @     �D@       @       @      �?     �C@      �?      L@              ?@      ,@      @      $@      @      @      �?      @      9@      @      5@              @      @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJH�SshG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK-hyh(h+K ��h-��R�(KK-��h��B�	                             �? �����?�           8�@                           @�`㖪�?y            �g@       
       	          033@�S�%3��?f            �c@                           �?l������?`            �b@                          �s@�t:ɨ�?T            �`@������������������������       �        J             ^@������������������������       ��q�q�?
             (@       	                     M@j���� �?             1@������������������������       �                      @������������������������       ��<ݚ�?             "@������������������������       �                     $@                           �O@ 	��p�?             =@������������������������       �                     7@                          �p@�q�q�?             @������������������������       �                     @������������������������       �                      @                            @:Vg{�?           �z@                          �a@`!'1��?�            �h@                           �?��s����?)            �O@                           �?�r����?            �F@������������������������       �X�<ݚ�?             "@������������������������       ��X�<ݺ?             B@                          `_@�q�q�?             2@������������������������       �                     @������������������������       �      �?	             (@              	          `ff@���y4F�?[            �`@                          `\@�חF�P�?T             _@������������������������       �b�2�tk�?             2@������������������������       ���-#���?I            �Z@                           �?�����H�?             "@������������������������       �                     @������������������������       �r�q��?             @!       &                   @[@�nq�o��?�            �l@"       #                     L@և���X�?	             ,@������������������������       �                     @$       %                    �?؇���X�?             @������������������������       �                     @������������������������       �                     �?'       *                    q@�n`���?�             k@(       )                   �d@r֛w���?d            `c@������������������������       �ܱ#_��?_            `b@������������������������       �                      @+       ,                    �?�g�y��?&             O@������������������������       �                     J@������������������������       �z�G�z�?             $@�t�bh�h(h+K ��h-��R�(KK-KK��ha�B�       Ps@      s@     �H@     `a@      6@      a@      (@      a@      @     �_@              ^@      @      @      @      $@               @      @       @      $@              ;@       @      7@              @       @      @                       @     @p@     �d@     �S@     @]@     �I@      (@     �C@      @      @      @      A@       @      (@      @      @              @      @      <@     @Z@      4@      Z@      &@      @      "@     @X@       @      �?      @              @      �?     �f@      I@      @       @              @      @      �?      @                      �?     �e@      E@     �\@      D@     �\@      @@               @      N@       @      J@               @       @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ�8�hG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK9hyh(h+K ��h-��R�(KK9��h��Bx                            Pb@���M#�?�           8�@                          �p@$��fF?�?�            @o@       
                    �?P�+���?n            �e@                           �?N֩	%��?3            @V@                           �?�GN�z�?             F@������������������������       �$��m��?             :@������������������������       ��X�<ݺ?             2@       	       	          `ff�?���X�K�?            �F@������������������������       �      �?             :@������������������������       �                     3@                          0b@�w>�
��?;            �T@                           [@8�Z$���?8            �S@������������������������       �                      @������������������������       ��?�'�@�?6             S@                           �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?                           �?ȵHPS!�?1            �S@                           �?�G�z��?             4@                          8s@z�G�z�?             $@������������������������       �                      @������������������������       �                      @                           t@�z�G��?             $@������������������������       �                     @������������������������       �                     @������������������������       �        %             M@       *                    @��>x7��?�            �v@       #                    �?�1����?�            `p@                            �? =[y��?}            �i@                          Xq@�����?.            �R@������������������������       �XB���?#             M@������������������������       �     ��?             0@!       "                    �? ����?O            @`@������������������������       �        '             P@������������������������       �Pa�	�?(            �P@$       '                   �_@^l��[B�?&             M@%       &                    �?��S���?	             .@������������������������       �                     @������������������������       �                      @(       )                    �?(L���?            �E@������������������������       �      �?             @������������������������       ��L���?            �B@+       2                    �?������?F            �Y@,       /                    �?R�}e�.�?%             J@-       .                    �?��.k���?             1@������������������������       �                      @������������������������       �                     "@0       1                    �K@؇���X�?            �A@������������������������       �X�Cc�?	             ,@������������������������       �                     5@3       6       
             �?�"U����?!            �I@4       5                    �P@r�q��?             8@������������������������       ��G��l��?             5@������������������������       �                     @7       8                    �?�<ݚ�?             ;@������������������������       �      �?             (@������������������������       �        
             .@�t�bh�h(h+K ��h-��R�(KK9KK��ha�B�       p@     `v@     @f@      R@     @[@     �O@      E@     �G@      $@      A@      "@      1@      �?      1@      @@      *@      *@      *@      3@             �P@      0@     �P@      (@               @     �P@      $@      �?      @              @      �?             @Q@      "@      &@      "@       @       @       @                       @      @      @              @      @              M@             �S@     �q@      6@      n@      "@     `h@      @     �P@       @      L@      @      &@       @      `@              P@       @      P@      *@     �F@      @       @      @                       @      @     �B@      @      @      @      A@     �L@      G@      C@      ,@       @      "@       @                      "@      >@      @      "@      @      5@              3@      @@      *@      &@      $@      &@      @              @      5@      @      @              .@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJUehG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK7hyh(h+K ��h-��R�(KK7��h��B                            Pb@&n.���?�           8�@              	          pff�?�<dۻC�?�             q@       
                    �?�H�a��?0            @U@                           @�X�<ݺ?!             K@                          �p@����?�?            �F@������������������������       �                    �D@������������������������       �      �?             @       	                    _@�<ݚ�?             "@������������������������       ��q�q�?             @������������������������       �                     @                          �Z@��a�n`�?             ?@������������������������       �                     @              	          833�?$�q-�?             :@������������������������       �        	             4@������������������������       ��q�q�?             @                          a@�����H�?v            �g@                           @,(��?K            �_@                           �?`2U0*��?I            @_@������������������������       ��LQ�1	�?             7@������������������������       ����J��?>            �Y@              	          `ff�?      �?              @������������������������       �                     �?������������������������       �                     �?                           �?j�g�y�?+             O@                           �?r�q��?             8@������������������������       �                     @������������������������       ��G�z��?             4@                           �?�KM�]�?             C@������������������������       �                     :@������������������������       ��q�q�?	             (@       *                    �L@���8S�?�            Pu@        '                   Ph@г����?�             o@!       $                    �?0������?�            @n@"       #       	          `ff@�t����?�            �i@������������������������       �,�8����?�            `i@������������������������       �                     �?%       &                    @P����?             C@������������������������       �                     2@������������������������       ���Q��?             4@(       )                    �?�q�q�?             @������������������������       �                      @������������������������       �                     @+       0                    @ܐ҆��??            @W@,       /       	          033@���3�E�?"             J@-       .                    �?�3Ea�$�?             G@������������������������       �l��\��?             A@������������������������       �      �?             (@������������������������       �                     @1       4                    �?���?            �D@2       3                   �`@$�q-�?             :@������������������������       �        
             ,@������������������������       �r�q��?             (@5       6                   �e@��S���?             .@������������������������       ��q�q�?	             (@������������������������       �                     @�t�bh�h(h+K ��h-��R�(KK7KK��ha�Bp       �q@     �t@     `h@     �S@      ;@      M@      @     �I@      �?      F@             �D@      �?      @       @      @       @      �?              @      8@      @              @      8@       @      4@              @       @      e@      5@     @^@      @      ^@      @      4@      @      Y@       @      �?      �?      �?                      �?     �G@      .@      *@      &@      @              "@      &@      A@      @      :@               @      @     �U@     �o@     �D@     �i@     �B@     �i@      8@     �f@      7@     �f@      �?              *@      9@              2@      *@      @      @       @               @      @              G@     �G@      .@     �B@      "@     �B@      @      ?@      @      @      @              ?@      $@      8@       @      ,@              $@       @      @       @      @       @      @        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ�)�rhG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK;hyh(h+K ��h-��R�(KK;��h��B�                             @&n.���?           8�@                           �?�(/���?�            Px@       
                    �?��\���?Q             a@                          Ps@4�B��?.            �R@              	          ���@��f/w�?(            �N@������������������������       �؇���X�?%             L@������������������������       �                     @       	                   �d@8�Z$���?             *@������������������������       ����Q��?             @������������������������       �                      @                          �Z@6uH���?#             O@                          �Y@      �?             @������������������������       �                     �?������������������������       �                     @                           �?XB���?              M@������������������������       �z�G�z�?             $@������������������������       �                     H@                           �?pe7����?�            �o@              	          033@�+$�jP�?>             [@                          �b@8�Z$���?;             Z@������������������������       ��^'�ë�?7            @X@������������������������       �؇���X�?             @������������������������       �                     @              	          hff @��Ή�ν?^             b@                           @��.N"Ҭ?Z            @a@������������������������       �`���i��?U            �`@������������������������       �r�q��?             @                           �?����X�?             @������������������������       �                      @������������������������       �                     @       ,                   �a@�ψX�F�?�            @l@        %                    [@��s�n�?D             Z@!       $                   �p@8�Z$���?
             *@"       #                    a@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     $@&       )                    �?x��B�R�?:            �V@'       (                    �?      �?	             0@������������������������       �                      @������������������������       �                     ,@*       +                     P@�}��L�?1            �R@������������������������       �        ,            �P@������������������������       �      �?              @-       4                    �?��C����?N            �^@.       1                   pb@Ɣ��Hr�?&            �M@/       0                   �^@�p ��?            �D@������������������������       �$��m��?             :@������������������������       �z�G�z�?	             .@2       3                    �?�����H�?             2@������������������������       �                     0@������������������������       �                      @5       8                   �_@Z���c��?(            �O@6       7                    �?      �?             0@������������������������       �                     @������������������������       �r�q��?	             (@9       :                    �?=QcG��?            �G@������������������������       �                     @@������������������������       �z�G�z�?	             .@�t�bh�h(h+K ��h-��R�(KK;KK��ha�B�       �q@     �t@     �[@     pq@     @T@     �K@      8@      I@      *@      H@       @      H@      @              &@       @      @       @       @             �L@      @      �?      @      �?                      @      L@       @       @       @      H@              =@      l@      4@      V@      0@      V@      $@     �U@      @      �?      @              "@      a@      @     �`@      @      `@      �?      @      @       @               @      @             �e@      K@     �X@      @      &@       @      �?       @               @      �?              $@              V@      @      ,@       @               @      ,@             �R@      �?     �P@              @      �?     @R@     �H@      7@      B@      5@      4@      "@      1@      (@      @       @      0@              0@       @              I@      *@      @      $@      @               @      $@      F@      @      @@              (@      @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJX"4qhG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK5hyh(h+K ��h-��R�(KK5��h��B�                             �?;�׊��?�           8�@                           @F�^Q��?�            ps@       
                    �?�G��l��?Y            `b@                           �?�q�q�?S            �`@              	          `ff@:�&���?4            �S@������������������������       ������H�?1             R@������������������������       �                     @       	       
             �?����|e�?             K@������������������������       ��<ݚ�?            �F@������������������������       ��q�q�?             "@������������������������       �                     .@                           �O@0��P�?e            �d@                          @[@hڛ�ʚ�?\            �b@                          0m@���Q��?             @������������������������       �                      @������������������������       �                     @                          �m@@��8��?Y             b@������������������������       �0G���ջ?!             J@������������������������       �        8             W@                          �^@�q�q�?	             .@              	          ����?z�G�z�?             @������������������������       �                     @������������������������       �                     �?                           �?ףp=
�?             $@������������������������       �z�G�z�?             @������������������������       �                     @       (                    �K@�I�w�"�?�             s@       !                   �a@      �?w             f@                           �?���!pc�?             6@������������������������       �                      @                           �^@և���X�?             ,@������������������������       �      �?              @������������������������       �                     @"       %                    @���j�?g            @c@#       $                    �?@�E�x�?b            `b@������������������������       �        '            �M@������������������������       ��zvܰ?;             V@&       '                   �j@����X�?             @������������������������       �                     @������������������������       ��q�q�?             @)       .       	          ����?     ��?L             `@*       +                    �?�q�q�?0            �S@������������������������       �                     "@,       -                    �L@�G�5��?-            @Q@������������������������       �p�ݯ��?
             3@������������������������       �ףp=
�?#             I@/       2                    @�z�G��?             I@0       1       	          ���@8�A�0��?             6@������������������������       �������?             1@������������������������       �                     @3       4       	          ���@@4և���?             <@������������������������       �                     :@������������������������       �                      @�t�bh�h(h+K ��h-��R�(KK5KK��ha�BP       �r@     �s@      l@     �U@     �Q@     @S@     �K@     @S@      ,@      P@       @      P@      @             �D@      *@     �A@      $@      @      @      .@             @c@      $@      b@      @      @       @               @      @             �a@      @     �H@      @      W@              $@      @      �?      @              @      �?              "@      �?      @      �?      @              R@      m@      &@     �d@      @      0@               @      @       @      @       @              @      @     �b@      @      b@             �M@      @     @U@       @      @              @       @      �?     �N@     �P@      :@      J@      "@              1@      J@      (@      @      @     �F@     �A@      .@      "@      *@      @      *@      @              :@       @      :@                       @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ;�3whG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK)hyh(h+K ��h-��R�(KK)��h��B�                	          ����?BM�e�x�?�           8�@                           �?t��g��?7           �~@       
       	          033�?V�a�� �?�            �s@                          Pb@���B���?�            �s@                          �\@^�JB=�?8            @T@������������������������       � �Cc}�?             <@������������������������       �~|z����?&            �J@       	                    �? ���?�            �l@������������������������       �`Ӹ����?4            �V@������������������������       �~F�̫�?X            �a@                          �\@؇���X�?             @������������������������       �                     �?������������������������       �                     @                           �?s8?U��?n            �e@                           `@*Mp����?C            �Y@������������������������       �                      @                           @��n%�4�?;            �W@������������������������       �      �?/             R@������������������������       �                     6@              	          ����?��oh���?+            @R@                          8p@b�2�tk�?             B@������������������������       �                     3@������������������������       �@�0�!��?             1@                          �_@@-�_ .�?            �B@������������������������       ��r����?
             .@������������������������       �                     6@       &                    @�C��2(�?O            @^@       !                    �F@�}�+r��?J            �\@                           �?���|���?             &@������������������������       �                      @                            @F@�<ݚ�?             "@������������������������       �                     @������������������������       �                      @"       %                    �?p� V�?B            �Y@#       $       
             �?z�G�z�?             $@������������������������       �                      @������������������������       �                      @������������������������       �        <            @W@'       (       
             �?����X�?             @������������������������       �                     @������������������������       �                      @�t�b��     h�h(h+K ��h-��R�(KK)KK��ha�B�       �p@     �u@     �c@      u@     �P@     �o@      N@     �o@      ?@      I@      @      9@      <@      9@      =@     @i@      @     �U@      9@      ]@      @      �?              �?      @              W@     �T@     �A@     �P@       @              ;@     �P@      ;@     �F@              6@     �L@      0@      6@      ,@      3@              @      ,@     �A@       @      *@       @      6@             �[@      &@      [@      @      @      @               @      @       @      @                       @     @Y@       @       @       @       @                       @     @W@               @      @              @       @        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ�3hG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK/hyh(h+K ��h-��R�(KK/��h��BH
                             @D^��#��?}           8�@                           �?�B7c�?�            �v@                           �?^����?            �E@                           �?X�Cc�?
             ,@������������������������       �                     "@������������������������       �                     @                           �?ܷ��?��?             =@������������������������       �                     2@	       
                    @I@���!pc�?             &@������������������������       �                      @������������������������       �                     @                          �[@tk~X��?�            @t@                           �E@�Q����?             D@������������������������       �                     @              
             �?���|���?            �@@������������������������       �d}h���?	             ,@������������������������       ��\��N��?             3@                           @K@�+�cP!�?�            �q@                          �`@h㱪��?c            �d@������������������������       �                     @������������������������       �@3����?a            @d@                          �c@�0�w�?P            �]@������������������������       ��n����?H            @Z@������������������������       �����X�?             ,@                            �?��K�[��?�             o@                          �p@ wVX(6�?`            @d@                           �?���c���?A             Z@������������������������       �        	             .@                          0a@4\�����?8            @V@������������������������       �d��0u��?'             N@������������������������       �XB���?             =@������������������������       �                     M@!       (                   pq@      �?5            �U@"       %                    @�萻/#�?+            �P@#       $                   �Z@��B����?#             J@������������������������       �                     @������������������������       ����Q��?             �F@&       '                    �?��S�ۿ?             .@������������������������       �                     (@������������������������       ��q�q�?             @)       ,       
             �?���y4F�?
             3@*       +                   e@@4և���?             ,@������������������������       �                     *@������������������������       �                     �?-       .                    �?���Q��?             @������������������������       �                      @������������������������       �                     @�t�bh�h(h+K ��h-��R�(KK/KK��ha�B�       �q@     �t@     �W@     q@      ?@      (@      @      "@              "@      @              :@      @      2@               @      @       @                      @     �O@     Pp@      5@      3@              @      5@      (@      &@      @      $@      "@      E@     @n@      @     �c@      @              @     �c@      B@     �T@      :@     �S@      $@      @     �g@     �L@     �b@      ,@     �V@      ,@      .@             �R@      ,@     �G@      *@      <@      �?      M@             �E@     �E@      <@     �C@      ;@      9@              @      ;@      2@      �?      ,@              (@      �?       @      .@      @      *@      �?      *@                      �?       @      @       @                      @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ� �NhG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK)hyh(h+K ��h-��R�(KK)��h��B�                             �?;�׊��?�           8�@                          0f@BSf���?�            r@       
                   Pb@|���~�?�             q@                           �?ܷ��?��?r            �e@                          �]@�c�Α�?             =@������������������������       �                     @������������������������       ����}<S�?             7@       	                    �? 	��p�?]             b@������������������������       ��>4և��?             <@������������������������       �@\�*��?H            @]@                           @�z�G��?D             Y@                           �M@      �?             E@������������������������       ��㙢�c�?             7@������������������������       ��KM�]�?             3@                           �L@Riv����?&             M@������������������������       ��ՙ/�?             5@������������������������       ��?�|�?            �B@������������������������       �        
             .@                           @vAƠB��?�            `t@              	          `ff@$%j����?�            �o@                           �?6uH���?�             o@                          �n@�q�q�?             .@������������������������       �r�q��?             (@������������������������       �                     @                          �d@`�q��־?�             m@������������������������       ��8'��?T            @^@������������������������       �        A             \@������������������������       �                     @       $       	          ����?b1<+�C�?/            @R@       !                   �a@�99lMt�?            �C@                           �`@z�G�z�?             $@������������������������       �                      @������������������������       �                      @"       #                   �f@V�a�� �?             =@������������������������       ��>4և��?             <@������������������������       �                     �?%       (                   H{@l��\��?             A@&       '                    �I@�FVQ&�?            �@@������������������������       �                     &@������������������������       ��C��2(�?             6@������������������������       �                     �?�t�bh�h(h+K ��h-��R�(KK)KK��ha�B�       �r@     �s@     @l@     �O@     @l@      H@     �c@      2@      5@       @              @      5@       @     �`@      $@      7@      @      \@      @     �Q@      >@      5@      5@      @      3@      1@       @     �H@      "@      *@       @      B@      �?              .@     �Q@      p@      9@     �l@      4@     �l@      @      $@       @      $@      @              .@     @k@      .@     �Z@              \@      @             �F@      <@      ,@      9@       @       @       @                       @      @      7@      @      7@      �?              ?@      @      ?@       @      &@              4@       @              �?�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ���bhG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK/hyh(h+K ��h-��R�(KK/��h��BH
                             �?��S���?�           8�@                           @&S��:�?�            �r@       
                    �?N�� ���?Q            �`@                          Ps@<�A+K&�?0             S@                           �?��IF�E�?)            �P@������������������������       ��'�`d�?            �@@������������������������       �                    �@@       	                    �N@���Q��?             $@������������������������       �؇���X�?             @������������������������       �                     @                           �?؇���X�?!             L@                           �?��S���?	             .@������������������������       ��n_Y�K�?             *@������������������������       �                      @������������������������       �                    �D@              	          ����?(�s���?m             e@                          �m@��<b���?             G@                           @G@     ��?
             0@������������������������       �                      @������������������������       �X�Cc�?	             ,@              	          ����?(;L]n�?             >@������������������������       �        
             2@������������������������       ��8��8��?             (@������������������������       �        R            �^@       (       	          033�?ld�@���?�            �s@       !                    �K@��W��?�            �q@                          �[@���1j	�?n            �e@                           �?�θ�?             :@������������������������       �                     @������������������������       ������?             3@                            c@��pBI�?^            @b@������������������������       �                     �?������������������������       �@��t��?]             b@"       %                    �?F��L�?F            @[@#       $                    �M@Du9iH��?            �E@������������������������       �      �?             @������������������������       �                    �C@&       '                   Po@�eP*L��?*            �P@������������������������       ��%^�?            �E@������������������������       ��㙢�c�?             7@)       .                    �?�������?             A@*       +                    �?���Q��?             .@������������������������       �                      @,       -                    b@��
ц��?
             *@������������������������       �      �?              @������������������������       �                     @������������������������       �        
             3@�t�bh�h(h+K ��h-��R�(KK/KK��ha�B�       �q@     �t@     `k@     @T@     �N@     �Q@      *@     �O@      @     �M@      @      :@             �@@      @      @      @      �?              @      H@       @      @       @      @       @       @             �D@             �c@      $@      B@      $@      @      "@       @              @      "@      =@      �?      2@              &@      �?     �^@              Q@     �n@     �E@     �m@      $@     @d@      @      4@              @      @      *@      @     �a@      �?              @     �a@     �@@      S@      @      D@      @      �?             �C@      >@      B@      &@      @@      3@      @      9@      "@      @      "@               @      @      @      @       @              @      3@        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ+�MhG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK9hyh(h+K ��h-��R�(KK9��h��Bx                             �?Pf�.���?�           8�@                           �?<���q�?�            0r@       
                    �?��J~��?W             b@                           b@fv�S��?2            �T@                           X@��n�?-            �R@������������������������       �                     @������������������������       �D��\��?+            �Q@       	                    �?����X�?             @������������������������       �r�q��?             @������������������������       �                     �?              	          ����?�? Da�?%            �O@                           @      �?             <@������������������������       ��z�G��?             $@������������������������       �        	             2@                          �Z@��?^�k�?            �A@������������������������       �                     �?������������������������       �                     A@                           �?�F��O�?_            @b@                           `@����D��?=            @W@                          �c@@-�_ .�?            �B@������������������������       �                     >@������������������������       �����X�?             @������������������������       �        %             L@                           @r�����?"            �J@                           �O@�q�q�?             @������������������������       �                      @������������������������       �                     @                          �b@��E�B��?            �G@������������������������       ��θ�?             :@������������������������       �                     5@       ,                    @tk~X��?�            @t@        %                   pc@��tM��?�            �o@!       $                    �N@�D��?B            �X@"       #                    �?�q�q�?1            �S@������������������������       ��G�5��?+            @Q@������������������������       �                     "@������������������������       �                     4@&       )       	          ����?@��z��?^            �c@'       (                   �d@���M�?4            @V@������������������������       ��	j*D�?	             *@������������������������       �P�Lt�<�?+             S@*       +                    @�\=lf�?*            �P@������������������������       �        &            �N@������������������������       �r�q��?             @-       2                    �?և���X�?2            �Q@.       /                   �`@��Q���?             D@������������������������       �                      @0       1       	          ����?�I�w�"�?             C@������������������������       �                     @������������������������       �     ��?             @@3       6                   �_@d��0u��?             >@4       5                   �a@j���� �?             1@������������������������       �                     @������������������������       ��C��2(�?             &@7       8                   �b@$�q-�?
             *@������������������������       ��q�q�?             @������������������������       �                     $@�t�bh�h(h+K ��h-��R�(KK9KK��ha�B�       �p@     �u@      j@     �T@     �R@     �Q@      3@     �O@      ,@     �N@      @              $@     �N@      @       @      @      �?              �?     �K@       @      5@      @      @      @      2@              A@      �?              �?      A@             �`@      (@     �V@       @     �A@       @      >@              @       @      L@             �E@      $@       @      @       @                      @     �D@      @      4@      @      5@             �O@     Pp@     �@@     �k@      :@      R@      :@      J@      1@      J@      "@                      4@      @     �b@      @     �T@      @      "@       @     �R@      �?     �P@             �N@      �?      @      >@      D@      &@      =@       @              "@      =@              @      "@      7@      3@      &@      @      $@      @              �?      $@      (@      �?       @      �?      $@        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJY]hG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK7hyh(h+K ��h-��R�(KK7��h��B                            pb@��O���?�           8�@                           �?�E��ӭ�?�             r@                          �c@4����?            �j@              	          pff�?      �?              @������������������������       �                      @������������������������       �                     @       
                    �?���x��?y            �i@       	                    @�w>�
��?-            �T@������������������������       �|��?���?             ;@������������������������       �h�����?             L@                          @[@ @|���?L            �^@������������������������       �      �?              @������������������������       �P�Lt�<�?F            �\@              	          `ff�?`�Q��?0            �R@                          Po@д>��C�?%             M@              	          pff�?������?            �D@������������������������       �                     :@������������������������       ��r����?	             .@                           �?��.k���?             1@������������������������       �z�G�z�?             @������������������������       ��q�q�?	             (@              	           33@@�0�!��?             1@                           �O@��S�ۿ?	             .@������������������������       �                     (@������������������������       ��q�q�?             @������������������������       �                      @       (                    �?������?�            pt@       #                    �?�2;�f�?D            �W@                           �c@Ȩ�I��?(            �J@                           �?�\��N��?             3@������������������������       �                     @������������������������       �r�q��?             (@!       "                   �d@�t����?             A@������������������������       �                     .@������������������������       ����y4F�?             3@$       '                    @���N8�?             E@%       &                   �c@8�Z$���?	             *@������������������������       ����Q��?             @������������������������       �                      @������������������������       �                     =@)       0       
             �?�'�f7��?�             m@*       -                    @^������?0            �Q@+       ,                    @L@R���Q�?             D@������������������������       �                     ?@������������������������       ��q�q�?             "@.       /       	          ����?���Q��?             >@������������������������       ����Q��?
             .@������������������������       �z�G�z�?             .@1       4                    �?�����H�?l            @d@2       3       	          ����?      �?C             X@������������������������       �����˵�?(            �M@������������������������       �                    �B@5       6                    �?�GN�z�?)            �P@������������������������       ��z�G��?             4@������������������������       ���<b�ƥ?             G@�t�bh�h(h+K ��h-��R�(KK7KK��ha�Bp        s@     ps@      j@      T@      g@      =@       @      @       @                      @     �f@      7@     �P@      0@      *@      ,@      K@       @     �\@      @      @      @     �[@      @      8@     �I@      $@      H@       @     �C@              :@       @      *@       @      "@      @      �?      @       @      ,@      @      ,@      �?      (@               @      �?               @      X@     �l@      K@     �D@      ,@     �C@      $@      "@              @      $@       @      @      >@              .@      @      .@      D@       @      &@       @      @       @       @              =@              E@     �g@      8@      G@      @      A@              ?@      @      @      2@      (@      @      "@      (@      @      2@      b@      @     @W@      @      L@             �B@      .@     �I@      ,@      @      �?     �F@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ4
hG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK7hyh(h+K ��h-��R�(KK7��h��B                            pb@�>$�*��?�           8�@                           �?�1��i�?�            �p@       
                   @\@t��eh��?t             g@                           �?��Zy�?            �C@                           �?      �?
             0@������������������������       �z�G�z�?             @������������������������       �                     &@       	       	          ���@8����?             7@������������������������       �        
             0@������������������������       �                     @              
             �?�F��O�?]            @b@              	          pff�?�FVQ&�?U            �`@������������������������       �8����?             7@������������������������       ���wڝ�?I            @[@              	          833�?����X�?             ,@������������������������       �                     @������������������������       ��C��2(�?             &@                          �a@������?6            @T@              	            �?T����1�?&             M@                           @HP�s��?             9@������������������������       �                     5@������������������������       �      �?             @                           �?�'�=z��?            �@@������������������������       �                     (@������������������������       ���s����?             5@                          0b@���}<S�?             7@������������������������       �        
             0@                           �?����X�?             @������������������������       ����Q��?             @������������������������       �                      @       *                    @&x�
�?�            �u@        %                    �?����y7�?�            @o@!       $                    �?P̏����?$            �L@"       #                   `\@D>�Q�?"             J@������������������������       ����Q��?             @������������������������       ���E�B��?            �G@������������������������       �                     @&       '                    @L@�-j'�?x             h@������������������������       �        Z             b@(       )                    �?�q�q�?             H@������������������������       ��G�z��?             4@������������������������       �h�����?             <@+       0                    �?:ɨ��?@            �X@,       /                    �O@4��?�?             J@-       .       	             �? "��u�?             I@������������������������       �     ��?             @@������������������������       �        
             2@������������������������       �                      @1       4                    i@JJ����?!            �G@2       3                    �?�����H�?             "@������������������������       �                     �?������������������������       �                      @5       6                    �?�s��:��?             C@������������������������       �     ��?             0@������������������������       �"pc�
�?             6@�t�bh�h(h+K ��h-��R�(KK7KK��ha�Bp       �p@     �u@      f@     @V@     �c@      =@      6@      1@      .@      �?      @      �?      &@              @      0@              0@      @             �`@      (@      _@       @      0@      @      [@      �?      $@      @              @      $@      �?      5@      N@      3@     �C@       @      7@              5@       @       @      1@      0@              (@      1@      @       @      5@              0@       @      @       @      @               @     @W@      p@      8@     @l@      ,@     �E@      "@     �E@      @       @      @     �D@      @              $@     �f@              b@      $@      C@      "@      &@      �?      ;@     @Q@      >@     �G@      @     �G@      @      =@      @      2@                       @      6@      9@      �?       @      �?                       @      5@      1@      @      *@      2@      @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ��;hG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK1hyh(h+K ��h-��R�(KK1��h��B�
                             �?BM�e�x�?           8�@                           �?2�t����?�            `q@       
                   �a@��S���?Q             ^@                           �?z�):���?@             Y@              	          ����?r٣����?(            �P@������������������������       �                     >@������������������������       �X�<ݚ�?             B@       	       	            �?�t����?             A@������������������������       �������?
             .@������������������������       �                     3@                           @ףp=
�?             4@                          pb@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     1@                          v@l{��b��?^            �c@                          �e@��}� �?\            `c@              	            �?P-�T6��?Y            �b@������������������������       �������?            �B@������������������������       �0�)AU��?C            �\@                          �g@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @       &                    �?tw>��<�?�            u@              	          `ff�?��n5V�?�            `k@                           �? 
��р�?i             e@                          �c@      �?e             d@������������������������       ���<�Ұ?^            `b@������������������������       ��n_Y�K�?             *@������������������������       �                     "@        #                    q@H%u��?$             I@!       "                   p@t��ճC�?             F@������������������������       �P���Q�?             D@������������������������       �      �?             @$       %                    �?      �?             @������������������������       �                     @������������������������       �                     @'       ,                    �K@:���W�?C            �]@(       +                   @e@�:pΈ��?             I@)       *                    h@8��8���?             H@������������������������       �X�<ݚ�?             "@������������������������       �                    �C@������������������������       �                      @-       0       	          `ff�?�������?'             Q@.       /                    �?ҳ�wY;�?            �I@������������������������       ����Q��?             >@������������������������       �                     5@������������������������       �        
             1@�t�bh�h(h+K ��h-��R�(KK1KK��ha�B       �p@     �u@     @j@      Q@      P@      L@      G@      K@      0@      I@              >@      0@      4@      >@      @      &@      @      3@              2@       @      �?       @      �?                       @      1@             @b@      (@     @b@      "@      b@      @     �@@      @      \@       @      �?      @              @      �?                      @      M@     pq@      0@     `i@      $@     �c@      $@     �b@      @     �a@      @       @              "@      @      F@      @     �D@       @      C@      �?      @      @      @              @      @              E@      S@      @     �E@      @     �E@      @      @             �C@       @             �A@     �@@      2@     �@@      2@      (@              5@      1@        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJS�)/hG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK5hyh(h+K ��h-��R�(KK5��h��B�                             �?�:�Ӛ��?�           8�@                           �?2��x[��?�            �x@                           �?`Pp�I�?�            �n@                           X@�ˡ�5��?*            �Q@������������������������       �                     @                           �D@�G�V�e�?(             Q@������������������������       �z�G�z�?             @������������������������       ��[|x��?$            �O@	                           q@<;n,��?w             f@
                          e@X�Հ�+�?[            �`@������������������������       ������?3            �R@������������������������       �        (            �N@                           �L@�p ��?            �D@������������������������       �                     8@������������������������       �ҳ�wY;�?             1@                           �?և���X�?^            `b@                           �?���� �?            �D@                           �?�G��l��?             5@������������������������       �������?             .@������������������������       �                     @������������������������       �                     4@                           �?���vq�?C            �Z@                           @`�q�0ܴ?            �G@������������������������       �                     C@������������������������       ��<ݚ�?             "@              	          033�?�ݜ����?%            �M@������������������������       �r�qG�?             H@������������������������       �                     &@       (                   �b@������?�            �k@       #       	          ����?�$�����?j            @d@       "                   �p@��:x���?>            �X@        !                   a@R=6�z�?$            @P@������������������������       �RB)��.�?            �E@������������������������       ��eP*L��?             6@������������������������       �                     A@$       '                    @ ������?,            �O@%       &                   `b@�nkK�?             7@������������������������       �                     6@������������������������       �                     �?������������������������       �                     D@)       .                    �?����*��?!            �M@*       -                   �d@�θ�?             :@+       ,                    �M@���N8�?             5@������������������������       �        	             2@������������������������       ��q�q�?             @������������������������       �                     @/       2                   `d@���|���?            �@@0       1                    �I@؇���X�?             5@������������������������       �      �?             @������������������������       �        	             1@3       4                   Pe@      �?             (@������������������������       �                      @������������������������       �      �?             @�t�bh�h(h+K ��h-��R�(KK5KK��ha�BP       `q@     u@     @[@     �q@      9@     �k@      (@     �M@      @              "@     �M@      @      �?      @      M@      *@     `d@      @      `@      @     �P@             �N@      @     �A@              8@      @      &@      U@     �O@      &@      >@      &@      $@      &@      @              @              4@     @R@     �@@     �F@       @      C@              @       @      <@      ?@      1@      ?@      &@              e@      J@     �a@      4@      T@      3@      G@      3@      A@      "@      (@      $@      A@              O@      �?      6@      �?      6@                      �?      D@              ;@      @@      @      4@      �?      4@              2@      �?       @      @              5@      (@      2@      @      �?      @      1@              @      "@               @      @      �?�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ[س=hG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK-hyh(h+K ��h-��R�(KK-��h��B�	                             �?r�a����?�           8�@                           �?f.i��n�?�            Py@                           �?�z����?�            @p@������������������������       �        <             Y@                          �_@��Q���?b             d@                          e@�r*e���?,            �R@������������������������       ��zv�X�?             F@������������������������       �                     >@	       
                   @`@�4���L�?6            �U@������������������������       �                     @������������������������       �\���(\�?2             T@                          �a@20J�Ws�?\             b@                           �?�KM�]�?             C@                          �`@      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                     >@                          �k@n�tl��?C            �Z@                           �?���?            �D@������������������������       �                     @������������������������       �(N:!���?            �A@                           �?4���C�?,            �P@������������������������       ���� ��?             ?@������������������������       �">�֕�?            �A@                            �?4?~�0��?�            @j@                           �?�X����?             F@                          �b@���y4F�?             C@������������������������       �                     7@                           �?��S���?
             .@������������������������       ����!pc�?             &@������������������������       �                     @������������������������       �                     @!       (                   �n@�/ C-��?l            �d@"       %                   �i@�w�"w��?2             S@#       $                   �\@@-�_ .�?            �B@������������������������       �z�G�z�?             $@������������������������       �                     ;@&       '                   �a@Hث3���?            �C@������������������������       ��θ�?             :@������������������������       �        	             *@)       ,                   �p@����?�?:            �V@*       +                   `]@���}<S�?             7@������������������������       �      �?             @������������������������       �                     3@������������������������       �        )            �P@�t�bh�h(h+K ��h-��R�(KK-KK��ha�B�       �r@     �s@     �_@     pq@      F@      k@              Y@      F@      ]@      ;@     �G@      ;@      1@              >@      1@     @Q@      @              &@     @Q@     �T@     �O@      A@      @      @      @              @      @              >@              H@     �M@      $@      ?@      @              @      ?@      C@      <@      ;@      @      &@      8@     �e@     �B@      >@      ,@      >@       @      7@              @       @      @       @      @                      @     �a@      7@     �K@      5@     �A@       @       @       @      ;@              4@      3@      4@      @              *@      V@       @      5@       @       @       @      3@             �P@        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJnխphG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK;hyh(h+K ��h-��R�(KK;��h��B�                             �?D^��#��?           8�@                           �?H��Ly��?�            �v@       
                    �?����&�?�            �p@                           �?���7M�?G            @]@              
             �?��
P��?            �A@������������������������       �      �?             0@������������������������       �p�ݯ��?             3@       	                    �?��1��?3            �T@������������������������       �                     :@������������������������       �����>4�?"             L@                          �c@�.(�i��?[            �b@                          k@f>�cQ�?(            �N@������������������������       �                     C@������������������������       ��û��|�?             7@                           @�E�����?3            �V@������������������������       �        +            �R@������������������������       ���S�ۿ?             .@                           �?~	~���?=            �X@                           �O@��t���?2            �S@                          �Z@������?-            �Q@������������������������       �                     �?������������������������       � ���g=�?,            @Q@                           @X�<ݚ�?             "@������������������������       �                     @������������������������       �                     @                          �`@�����?             3@������������������������       �                     @                          �f@�r����?	             .@������������������������       �                     *@������������������������       �                      @       .       	          033�?\�DD��?�             o@        '                    �?��J�fj�?I            �[@!       $                   @[@�I�w�"�?             C@"       #                    �?r�q��?             @������������������������       �                     �?������������������������       �                     @%       &                   �Z@      �?             @@������������������������       �                      @������������������������       ���S�ۿ?             >@(       +                   �b@p�}�ޤ�?,            @R@)       *                    �?���Q��?             .@������������������������       �                     @������������������������       �"pc�
�?             &@,       -                    �?д>��C�?              M@������������������������       ��eP*L��?             6@������������������������       �                     B@/       6                    @D��*�4�?W            @a@0       3                    @J@z�G�z�?            �F@1       2                    �?r�q��?             @������������������������       �                     @������������������������       �                     �?4       5                   �r@��-�=��?            �C@������������������������       �г�wY;�?             A@������������������������       ����Q��?             @7       8                    �?�L��ȕ?<            @W@������������������������       �        1             S@9       :                     N@�IєX�?             1@������������������������       �                     (@������������������������       �z�G�z�?             @�t�bh�h(h+K ��h-��R�(KK;KK��ha�B�       �q@     �t@     @[@     p@      C@     �l@      <@     @V@      1@      2@      $@      @      @      (@      &@     �Q@              :@      &@     �F@      $@     �a@      "@      J@              C@      "@      ,@      �?     @V@             �R@      �?      ,@     �Q@      ;@     @P@      ,@     �N@      "@              �?     �N@       @      @      @              @      @              @      *@      @               @      *@              *@       @              f@     @R@      H@     �O@      =@      "@      �?      @      �?                      @      <@      @               @      <@       @      3@      K@      "@      @              @      "@       @      $@      H@      $@      (@              B@      `@      $@      B@      "@      �?      @              @      �?             �A@      @     �@@      �?       @      @      W@      �?      S@              0@      �?      (@              @      �?�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ�[�.hG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK/hyh(h+K ��h-��R�(KK/��h��BH
                             @�85�r��?�           8�@                           �?*��&��?�            `w@       
       	          ���@D��\��?�            �q@                           @L@�fɠ��?�            �p@                          �`@P����?p             f@������������������������       �      �?              @������������������������       �@�����?j             e@       	                    q@��+7��?>             W@������������������������       �d�;lr�?*            �O@������������������������       �П[;U��?             =@              
             �?�r����?	             .@                           �G@����X�?             @������������������������       �                     �?������������������������       �r�q��?             @������������������������       �                      @                          �Z@���X�K�?7            �V@                           �?�q�q�?             @              	          033�?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @                           �?0,Tg��?3             U@                           �?��hJ,�?)             Q@������������������������       �������?            �D@������������������������       ��<ݚ�?             ;@                           �?      �?
             0@������������������������       �                     "@������������������������       �և���X�?             @       &       	          pff�? -B��j�?�             n@                          �a@��j��?/            @S@������������������������       �                      @        #                    �?bKv���?*            @Q@!       "                    @L@�xGZ���?            �A@������������������������       �������?             1@������������������������       ��q�q�?	             2@$       %                   �b@H�V�e��?             A@������������������������       ��z�G��?             $@������������������������       �                     8@'       (                   �l@ĴF���?f            �d@������������������������       �        &             Q@)       ,                    �N@8��8���?@             X@*       +                   pm@����1�?1            @R@������������������������       ��q�q�?             @������������������������       ������?-            �P@-       .                   �]@8����?             7@������������������������       �                     @������������������������       �z�G�z�?             4@�t�bh�h(h+K ��h-��R�(KK/KK��ha�B�       �r@     �s@      Z@     �p@      D@     �n@      ;@     @n@      @     �e@       @      @      �?      e@      8@      Q@      &@      J@      *@      0@      *@       @      @       @              �?      @      �?       @              P@      :@       @      @       @       @       @                       @               @      O@      6@      M@      $@     �B@      @      5@      @      @      (@              "@      @      @      h@      H@     �E@      A@               @     �E@      :@      0@      3@      @      *@      (@      @      ;@      @      @      @      8@             �b@      ,@      Q@             �T@      ,@     �P@      @       @      @      P@      @      0@      @              @      0@      @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ��=hG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK1hyh(h+K ��h-��R�(KK1��h��B�
                             �?D^��#��?y           8�@                          pb@�0�~��?�             v@              	          pff�?���� �?J             _@                           �?     ��?             H@                           �K@�X���?             F@������������������������       �                     1@������������������������       �X�<ݚ�?             ;@������������������������       �                     @	                           @>A�F<�?/             S@
                            L@
j*D>�?             :@������������������������       ��r����?             .@������������������������       �"pc�
�?             &@              	          `ff@ "��u�?             I@������������������������       �                    �E@������������������������       �և���X�?             @                           @�?�'�@�?�            �l@                           �M@�f����?v             g@              	          033�?��X8��?c            @c@������������������������       �@�`%���?_            `b@������������������������       �����X�?             @                          �a@�4�����?             ?@������������������������       ��\��N��?             3@������������������������       �                     (@                          �p@�&!��?            �E@              
             �?�<ݚ�?             ;@������������������������       �      �?	             (@������������������������       �                     .@                           �?     ��?	             0@������������������������       ��eP*L��?             &@������������������������       �                     @       *       
             �?�ը��?�            pp@        %                    �?�r����?b            �d@!       "                    �O@����˵�?J            �]@������������������������       �        <            �W@#       $                    �?      �?             8@������������������������       ��q�q�?             @������������������������       ������H�?             2@&       '                    �?"Ae���?            �G@������������������������       �                     @(       )                    @R���Q�?             D@������������������������       �4?,R��?             B@������������������������       �                     @+       0                    @X�Cc�?:            �X@,       /                    �P@�q�q�?4             U@-       .                    �?      �?+            �Q@������������������������       �H�V�e��?             A@������������������������       ��<ݚ�?             B@������������������������       �        	             ,@������������������������       �                     ,@�t�bh�h(h+K ��h-��R�(KK1KK��ha�B       �q@     �t@     �Z@     �n@     @S@     �G@      .@     �@@      .@      =@              1@      .@      (@              @      O@      ,@      .@      &@      *@       @       @      "@     �G@      @     �E@              @      @      >@     �h@      *@     �e@      @     �b@      �?     @b@       @      @      $@      5@      $@      "@              (@      1@      :@      @      5@      @      @              .@      &@      @      @      @      @             @f@     @U@     �a@      6@      \@      @     �W@              2@      @       @      @      0@       @      ?@      0@              @      ?@      "@      ?@      @              @     �A@     �O@     �A@     �H@     �A@     �A@      ;@      @       @      <@              ,@              ,@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ��(hG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK5hyh(h+K ��h-��R�(KK5��h��B�                             �?JGC8{��?�           8�@                          �b@,�ѳ�?�             q@                           �?p`q�q��?e            �c@                          `c@h�����?E             \@������������������������       �        9            @V@              	          `ff�?�㙢�c�?             7@������������������������       �                     $@������������������������       ��	j*D�?             *@	              	          ����?�û��|�?              G@
                          �b@R�}e�.�?             :@������������������������       ���2(&�?             6@������������������������       �                     @              	          033�?�G�z��?             4@������������������������       �r�q��?	             (@������������������������       �      �?              @                          �p@p9W��S�?O            �\@                           @؇���X�?-            �O@                           n@���C��?%            �J@������������������������       �b�h�d.�?            �A@������������������������       �                     2@                           d@�z�G��?             $@������������������������       �؇���X�?             @������������������������       ��q�q�?             @                           �?��.k���?"            �I@                          @r@�lg����?            �E@������������������������       ��d�����?             3@������������������������       ��8��8��?             8@������������������������       �                      @       (                    �?3��9�?�            pu@       %                    f@v���6h�?�            `j@       "                    �?@�0�!��?�            �i@        !                    @������?j            �d@������������������������       ��Z]]Y�?X            �`@������������������������       ��z�G��?             >@#       $                    @      �?             D@������������������������       �X�Cc�?             <@������������������������       �r�q��?             (@&       '                    �M@؇���X�?             @������������������������       �                     @������������������������       �                     �?)       0                    �?�N2�,��?O            �`@*       -                    �O@r�q��?)            �S@+       ,                   @[@���N8�?             �O@������������������������       �      �?             @������������������������       �                    �L@.       /                    @P@�q�q�?	             .@������������������������       �                     @������������������������       �      �?             $@1       4       	          033�?������?&             K@2       3                    @Du9iH��?            �E@������������������������       ��?�|�?            �B@������������������������       ��q�q�?             @������������������������       �                     &@�t�bh�h(h+K ��h-��R�(KK5KK��ha�BP       �q@     �t@     �c@     @\@     �_@      @@      [@      @     @V@              3@      @      $@              "@      @      2@      <@      @      3@      @      3@      @              &@      "@      $@       @      �?      @     �@@     @T@      "@      K@      @     �G@      @      =@              2@      @      @      �?      @       @      �?      8@      ;@      0@      ;@      ,@      @       @      6@       @             @^@     �k@      E@      e@      B@      e@      0@     �b@      @     �_@      "@      5@      4@      4@      $@      2@      $@       @      @      �?      @                      �?     �S@     �J@     @P@      *@      N@      @      @      @     �L@              @      $@              @      @      @      ,@      D@      @      D@      �?      B@       @      @      &@        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ���~hG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK3hyh(h+K ��h-��R�(KK3��h��B(                            Pb@��>�'��?�           8�@                           �?��]��9�?�            pp@                           @X�<ݚ�?A            �X@                           @H@�'N��?(            �N@������������������������       �                     1@                            P@�zv�X�?             F@������������������������       ��X����?             6@������������������������       ��C��2(�?             6@	       
                    �L@p9W��S�?             C@������������������������       �        	             ,@              	          hff�?r�q��?             8@������������������������       �                     @������������������������       �������?             1@                           �?������?d            �d@                           `@��K˱F�?X            �a@                          �_@����p�?)             Q@������������������������       �        "             K@������������������������       �X�Cc�?             ,@������������������������       �        /            �R@                           �?�G��l��?             5@                          �`@X�Cc�?             ,@������������������������       �                     @������������������������       �                     "@                           �?����X�?             @������������������������       �                     �?������������������������       �r�q��?             @       *                    �?�GN��?�             v@       #                    �?j(���?�            @s@                           0n@��}����?6            �X@              	          `ff@�r����?            �F@������������������������       ��ʈD��?            �E@������������������������       �                      @!       "                   `u@|��?���?             K@������������������������       ��û��|�?             G@������������������������       �                      @$       '                   �l@T�fU���?�             j@%       &                    �?�ȉo(��?;            �V@������������������������       �r�q��?             8@������������������������       �        ,            �P@(       )                   �d@F�4�Dj�?T            �]@������������������������       �4Ky\�?O            @\@������������������������       �                     @+       2                   �o@���!pc�?             F@,       /                    @
;&����?             7@-       .                   �d@z�G�z�?             $@������������������������       �                      @������������������������       �                      @0       1                    @�	j*D�?             *@������������������������       �                     "@������������������������       �                     @������������������������       �                     5@�t�bh�h(h+K ��h-��R�(KK3KK��ha�B0       �q@     �t@      h@     �Q@      F@     �K@      1@      F@              1@      1@      ;@      .@      @       @      4@      ;@      &@      ,@              *@      &@              @      *@      @     �b@      0@     @a@      @     �O@      @      K@              "@      @     �R@              $@      &@      @      "@      @                      "@      @       @              �?      @      �?      W@     @p@      N@      o@      A@     @P@      @     �C@      @     �C@       @              <@      :@      <@      2@               @      :@     �f@      @     �U@      @      4@             �P@      6@      X@      1@      X@      @              @@      (@      &@      (@       @       @       @                       @      "@      @      "@                      @      5@        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJCLUhG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK1hyh(h+K ��h-��R�(KK1��h��B�
                            �a@��a��?�           8�@              	          ����?�1{�Z(�?�            @i@       
                    �P@<W#.m��?C            @Z@                           �?���!���?=            �W@                           @\�����?%            �K@������������������������       �ڡR����?!            �H@������������������������       �                     @       	                    @8�Z$���?            �C@������������������������       � >�֕�?            �A@������������������������       �                     @������������������������       �                     &@                           @h�a��?@            @X@                           �?д>��C�?             =@                           �?�q�q�?             @������������������������       �                     @������������������������       �                      @                           �?�nkK�?             7@������������������������       ��q�q�?             @������������������������       �                     4@������������������������       �        ,             Q@       $                    @"7r�@��?�            �y@                           �?    �/�?�             p@              	          033@Z��Yo��?*             O@                           �?R�}e�.�?$             J@������������������������       �z�G�z�?             D@������������������������       ��q�q�?	             (@                           @F@ףp=
�?             $@������������������������       �                     @������������������������       �z�G�z�?             @       !                   �d@������?x            @h@                           �b@P�#�Z�?>            �Y@������������������������       �ܷ��?��?             =@������������������������       ��1��u�?-            @R@"       #                   �_@�����?:             W@������������������������       �                     H@������������������������       �`���i��?             F@%       ,                   xq@�(T���?[            �c@&       )                    �?��C����?H            �^@'       (                    �?(2��R�?!            �M@������������������������       �      �?             0@������������������������       � �#�Ѵ�?            �E@*       +       	          ����?b����?'            �O@������������������������       ��t����?             A@������������������������       �����"�?             =@-       0                    @K@(N:!���?            �A@.       /                    �?�q�q�?             (@������������������������       �                      @������������������������       ����Q��?             $@������������������������       �                     7@�t�bh�h(h+K ��h-��R�(KK1KK��ha�B       �r@     �s@     �b@     �I@     �M@      G@     �M@     �A@      :@      =@      4@      =@      @             �@@      @     �@@       @              @              &@      W@      @      8@      @       @      @              @       @              6@      �?       @      �?      4@              Q@             �b@     `p@     �G@      j@      7@     �C@      ,@      C@      @     �@@      @      @      "@      �?      @              @      �?      8@     @e@      7@     �S@      @      :@      4@     �J@      �?     �V@              H@      �?     �E@      Z@     �J@     @R@     �H@     �I@       @      $@      @     �D@       @      6@     �D@      @      >@      2@      &@      ?@      @       @      @       @              @      @      7@        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ���hG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK5hyh(h+K ��h-��R�(KK5��h��B�                
             �?���i��?           8�@                          Pb@���v�?�            @t@              	          pff�?bۘ�W^�?�            @j@                           �?ڡR����?            �H@������������������������       �        
             0@                           @<���D�?            �@@������������������������       �                     9@������������������������       �      �?              @	                           �Q@���}<S�?k             d@
                           @��e3���?i            �c@������������������������       �D>�Q�?#             J@������������������������       ��O4R���?F            �Z@������������������������       �                     @                           @A�b��?G            �\@                           �?~X�<��?*             R@                           �?8�A�0��?             6@������������������������       ��	j*D�?             *@������������������������       �                     "@                          0g@z�G�z�?             I@������������������������       ��z�G��?             $@������������������������       ���(\���?             D@                          �p@�q�q�?             E@                          �c@���>4��?             <@������������������������       �b�2�tk�?             2@������������������������       �z�G�z�?             $@                          �]@@4և���?	             ,@������������������������       �                     �?������������������������       �                     *@       (                    �?�q4���?�            0r@       %                    �?��j2��?<            @Y@       "                   Hq@f1r��g�?#            �J@        !                   �[@ qP��B�?            �E@������������������������       ������H�?             "@������������������������       �                     A@#       $                    @O@�z�G��?             $@������������������������       �      �?              @������������������������       �                      @&       '                    �?      �?             H@������������������������       �                     @������������������������       �                     E@)       .                    @�¦�{��?v            �g@*       +                    @G@8$�s���?g            `d@������������������������       �                    �I@,       -                   �c@��X��?H             \@������������������������       �                     �?������������������������       ����l��?G            �[@/       2                   @b@�q�q�?             ;@0       1                   �`@�q�q�?             (@������������������������       �                     @������������������������       �                     @3       4                   �q@�r����?             .@������������������������       �@4և���?
             ,@������������������������       �                     �?�t�bh�h(h+K ��h-��R�(KK5KK��ha�BP       0r@     @t@     �k@     @Y@      f@      A@      =@      4@              0@      =@      @      9@              @      @     `b@      ,@     `b@      &@     �E@      "@      Z@       @              @     �G@     �P@      3@     �J@      "@      *@      "@      @              "@      $@      D@      @      @      @     �B@      <@      ,@      .@      *@      @      &@       @       @      *@      �?              �?      *@              Q@     �k@      I@     �I@       @     �F@      �?      E@      �?       @              A@      @      @      @      �?               @      E@      @              @      E@              2@     �e@      "@     @c@             �I@      "@     �Y@      �?               @     �Y@      "@      2@      @      @      @                      @       @      *@      �?      *@      �?        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ"�a,hG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK9hyh(h+K ��h-��R�(KK9��h��Bx                             �?��O���?�           8�@              	          pff�?��Ӊ�?�            �r@       
                    @xO�a���?J            @[@                          `a@p�ݯ��?)            �L@                          �Z@��Q��?             4@������������������������       �                     @������������������������       �     ��?
             0@       	                    �?���@��?            �B@������������������������       ��}�+r��?             3@������������������������       �b�2�tk�?             2@                           �?θ	j*�?!             J@                          �m@      �?             6@������������������������       �8�Z$���?             *@������������������������       �                     "@                          8p@z�G�z�?             >@������������������������       ��}�+r��?             3@������������������������       ��eP*L��?             &@                           �?,���$�?z            @h@                           �C@r�����?            �J@������������������������       �                     @                          �_@�q��/��?            �H@������������������������       �      �?              @������������������������       ���p\�?            �D@                           f@�lm�9�?]            �a@                           �E@ aqk+�?\            `a@������������������������       ��C��2(�?             &@������������������������       �     ��?V             `@������������������������       �                      @       ,                    @���5��?�            �s@       %                    �?x���� �?�             n@       "                   �d@f��>���?:            @U@        !       	          `ff�?L
�q��?(            �M@������������������������       ���|�5��?             �G@������������������������       �      �?             (@#       $                    �K@ ��WV�?             :@������������������������       �                     5@������������������������       �z�G�z�?             @&       )                    �?(�����?b            `c@'       (                   �`@և���X�?             @������������������������       �                     @������������������������       �                     @*       +                   Pd@,N�_� �?^            �b@������������������������       ��k�'7��?'            �L@������������������������       �        7            �V@-       2                    b@)O���?0             R@.       /                   @[@�û��|�?             G@������������������������       �                     @0       1                   �a@�(�Tw��?            �C@������������������������       �        
             1@������������������������       �      �?             6@3       6                    �?�θ�?             :@4       5                   c@z�G�z�?             4@������������������������       ��q�q�?             @������������������������       �        
             ,@7       8                   `c@�q�q�?             @������������������������       �                     @������������������������       �                      @�t�b���      h�h(h+K ��h-��R�(KK9KK��ha�B�        s@     ps@     �m@     �P@      L@     �J@      5@      B@      *@      @              @      *@      @       @      =@      �?      2@      @      &@     �A@      1@      &@      &@       @      &@      "@              8@      @      2@      �?      @      @     �f@      ,@     �E@      $@              @     �E@      @      @      @      C@      @      a@      @      a@       @      $@      �?     �_@      �?               @      Q@     �n@      A@     �i@      5@      P@      4@     �C@      &@      B@      "@      @      �?      9@              5@      �?      @      *@     �a@      @      @              @      @              $@     @a@      $@     �G@             �V@      A@      C@      <@      2@              @      <@      &@      1@              &@      &@      @      4@      @      0@      @       @              ,@       @      @              @       @        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ�8�hhG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK1hyh(h+K ��h-��R�(KK1��h��B�
                             @K@r�a����?�           8�@                           @��?����?�            `r@                           �?x�x
.L�?            �i@                           �?p�ݯ��?&            �L@������������������������       �                     5@                           �?�q�q�?             B@������������������������       ����|���?             6@������������������������       �@4և���?	             ,@	                           c@ �ޫ��?Y            �b@
                           @G@      �?              @������������������������       �                     �?������������������������       �                     �?                          c@@�E�x�?W            `b@������������������������       ��8��8��?             B@������������������������       �        B            �[@                          0b@�������?=             V@                           �I@�?�|�?            �B@������������������������       �                     <@                           �?�����H�?             "@������������������������       �                     �?������������������������       �                      @                          @[@�q�q�?#            �I@������������������������       �                     @                           �?�GN�z�?             F@������������������������       �J�8���?             =@������������������������       �                     .@       (                    �?r�0?��?�            t@       !                    @�#}���?y            �g@                            @�z�G��?L             ^@                           �?����՟�?F            @[@������������������������       ��eP*L��?             &@������������������������       ��[$�G�?A            �X@������������������������       �                     &@"       %                    @�ګH9�?-            �Q@#       $                   �a@z�G�z�?(            @P@������������������������       �v�X��?             F@������������������������       �                     5@&       '       	          ����?r�q��?             @������������������������       �                     �?������������������������       �                     @)       0                    @ȵHPS!�?N            @`@*       -       	          ����?R�xE��?M            �_@+       ,                   �_@\X��t�?             7@������������������������       �                      @������������������������       ��q�q�?             .@.       /                   v@ pƵHP�?>             Z@������������������������       ��K}��?<            �Y@������������������������       �      �?              @������������������������       �                     @�t�bh�h(h+K ��h-��R�(KK1KK��ha�B       �r@     �s@     �W@     �h@      9@     �f@      5@      B@              5@      5@      .@       @      ,@      *@      �?      @      b@      �?      �?              �?      �?              @      b@      @     �@@             �[@     �Q@      2@      B@      �?      <@               @      �?              �?       @              A@      1@              @      A@      $@      3@      $@      .@             �i@     @]@     @V@     �Y@      B@      U@      9@      U@      @      @      3@     �S@      &@             �J@      2@      J@      *@      ?@      *@      5@              �?      @      �?                      @     �\@      .@     �\@      (@      *@      $@       @              @      $@     �Y@       @     @Y@      �?      �?      �?              @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJP�dhG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK/hyh(h+K ��h-��R�(KK/��h��BH
                             �?��>�'��?           8�@              	          033�?x%[VY[�?�            �x@       
                    �?z�G�z�?�            0v@                           @����X��?�            �n@                          xt@P�2E��?{            `h@������������������������       ��˫���?s             g@������������������������       ����|���?             &@       	                     I@�"U����?            �I@������������������������       ��q�q�?             5@������������������������       �r�q��?             >@                           �?͍�@��?D            @[@                          �`@�θ�?"             J@������������������������       �                     (@������������������������       ��z�G��?             D@                          �l@�}�+r��?"            �L@������������������������       �     ��?
             0@������������������������       �                    �D@              	          `ff@v�X��?             F@                           �E@���y4F�?             C@������������������������       �                      @              
             �?r�q��?             B@������������������������       �      �?             @������������������������       �ףp=
�?             >@                           �?r�q��?             @������������������������       �                     @������������������������       �                     �?       &       	            �?BMĹ��?�             k@       !                   �b@��.k���?#            �I@              	          833�?��2(&�?             6@������������������������       �        
             (@                           �\@�z�G��?             $@������������������������       �                     @������������������������       �                     @"       #                    �?�c�Α�?             =@������������������������       �                     (@$       %                   `[@��.k���?             1@������������������������       �                     @������������������������       �և���X�?             ,@'       *                   �Z@�FVQ&�?d            �d@(       )                    �M@և���X�?             @������������������������       �                     @������������������������       �                     @+       .                    @��o;���?_            �c@,       -       
             �? ���l��?\            `c@������������������������       �`����֜?S            �a@������������������������       ��r����?	             .@������������������������       �                     @�t�bh�h(h+K ��h-��R�(KK/KK��ha�B�       �q@     �t@     �Y@     �r@     �Q@     �q@      <@     @k@      "@     @g@      @     `f@      @      @      3@      @@      ,@      @      @      9@     �E@     �P@      D@      (@      (@              <@      (@      @      K@      @      *@             �D@      ?@      *@      >@       @               @      >@      @      @      @      ;@      @      �?      @              @      �?             �f@      A@      ;@      8@      3@      @      (@              @      @              @      @               @      5@              (@       @      "@              @       @      @     `c@      $@      @      @              @      @             �b@      @     �b@      @     @a@       @      *@       @              @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ�g?BhG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK1hyh(h+K ��h-��R�(KK1��h��B�
                             @�:�Ӛ��?�           8�@                           �?Zfc��?�            x@                           �?     8�?X             `@                           �?P����?             C@              	          033�?<ݚ)�?             B@������������������������       ���a�n`�?             ?@������������������������       �z�G�z�?             @������������������������       �                      @	                           �?$�ݏ^��?9            �V@
                          �f@��V#�?            �E@������������������������       �                     @������������������������       ����@��?            �B@������������������������       �                    �G@                           �K@h�L�2��?�            p@                           c@0�)AU��?e            `e@������������������������       �                      @                          c@@�����?d             e@������������������������       �P�Lt�<�?             C@������������������������       �        O            ``@                           �?��|\�d�?4            �U@                          @b@�����H�?             "@������������������������       �                      @������������������������       �                     �?                          �p@��مD�?/            @S@������������������������       ��q��/��?            �H@������������������������       ���>4և�?             <@       *       	          033�?���?�            �l@       #                    �?Zz�����?;            @U@                            �K@f.i��n�?             �F@                          �p@��2(&�?             6@������������������������       �        
             .@������������������������       �և���X�?             @!       "       	          pff�?
;&����?             7@������������������������       �����X�?	             ,@������������������������       ������H�?             "@$       '                   �l@�z�G��?             D@%       &                    �?�θ�?	             *@������������������������       �                     @������������������������       �                     $@(       )                    �N@�>����?             ;@������������������������       � �q�q�?             8@������������������������       ��q�q�?             @+       ,                    �?�������?]             b@������������������������       �        G            �\@-       .                    @I@d��0u��?             >@������������������������       �                     @/       0                   �l@r�q��?             8@������������������������       �                      @������������������������       �     ��?             0@�t�bh�h(h+K ��h-��R�(KK1KK��ha�B       `q@     u@     �Y@     �q@     �R@      K@      *@      9@      &@      9@      @      8@      @      �?       @             �N@      =@      ,@      =@      @               @      =@     �G@              <@     �l@      @      e@       @              �?      e@      �?     �B@             ``@      9@     �N@       @      �?       @                      �?      1@      N@      @     �E@      &@      1@      f@      K@      E@     �E@      ,@      ?@      @      3@              .@      @      @      &@      (@      $@      @      �?       @      <@      (@      @      $@      @                      $@      9@       @      7@      �?       @      �?     �`@      &@     �\@              3@      &@      @              *@      &@       @              @      &@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ1�.hG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK1hyh(h+K ��h-��R�(KK1��h��B�
                             �?���i��?�           8�@       	                    �?^Z�sl�?�            �r@                          hs@X)0���?V            �`@                           �?�p ��?O            �^@                           �?��J�fj�?J            �[@������������������������       ���.��?-            �N@������������������������       ��+e�X�?             I@������������������������       �                     (@������������������������       �                     &@
                          pb@\�>���?n            �d@              
             �?X�Հ�+�?\            �`@                          �Z@ ,V�ނ�?U            �_@������������������������       ����N8�?             5@������������������������       �        H            @Z@                          �a@�<ݚ�?             "@������������������������       �                     @������������������������       ��q�q�?             @                           �?���@M^�?             ?@                          @`@���Q��?             4@������������������������       �      �?              @������������������������       �      �?	             (@������������������������       �                     &@       $                   �k@<-{)��?�            �s@                           �?�?�P�a�?I             ^@                          0g@��S�ۿ?5            �V@              	          hff@r�q��?             >@������������������������       �                     9@������������������������       �                     @                          �b@ �.�?Ƞ?&             N@������������������������       �        #            �L@������������������������       ��q�q�?             @        #                    �?������?             >@!       "       	          833�?H%u��?             9@������������������������       �                     5@������������������������       �      �?             @������������������������       �                     @%       *                    �K@Z��:��?{            `h@&       )                   �e@L紂P�?=            �Y@'       (       	          ���@ i���t�?;            �X@������������������������       � rpa�?8            @W@������������������������       �                     @������������������������       �                     @+       .                   �d@�g�y��?>            @W@,       -       	          033�?�W����?5            �T@������������������������       ��Ƀ aA�?'            �M@������������������������       ���<b���?             7@/       0                    �?"pc�
�?	             &@������������������������       �                     "@������������������������       �                      @�t�bh�h(h+K ��h-��R�(KK1KK��ha�B       0r@     @t@     @k@     �T@     �Q@     �O@      N@     �O@      H@     �O@      $@     �I@      C@      (@      (@              &@             `b@      3@      `@      @     @^@      @      0@      @     @Z@              @       @      @              �?       @      3@      (@       @      (@      @      @      @      "@      &@             @R@     @n@      ,@     �Z@      @      U@      @      9@              9@      @              �?     �M@             �L@      �?       @       @      6@      @      6@              5@      @      �?      @             �M@      a@      ,@      V@      $@      V@      @      V@      @              @             �F@      H@     �E@     �C@      9@      A@      2@      @       @      "@              "@       @        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJg�)hG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK1hyh(h+K ��h-��R�(KK1��h��B�
                
             �?|��z��?�           8�@              	          033�?"�a�5M�?�            t@                           @��V�I��?;            �W@                          @]@�q�q�?&            �L@������������������������       �                     *@                           �K@��2(&�?             F@������������������������       �                    �@@������������������������       ��eP*L��?
             &@	                           �?؀�:M�?            �B@
                           �?���B���?             :@������������������������       ����N8�?             5@������������������������       �                     @                          �n@"pc�
�?             &@������������������������       �                     @������������������������       ����Q��?             @                           �Q@�>:���?�            `l@                           @��G���?�            �k@              	          `ff @�O�w���?8            �V@������������������������       �6C�z��?$            �L@������������������������       ���hJ,�?             A@                          h~@�-�[�?T            ``@������������������������       � �#�Ѵ�?S             `@������������������������       �                      @������������������������       �                     @       &                    �?���c�H�?�            `r@                           @X�<ݚ�?<            �V@              	          ����?�GN�z�?             F@                            P@����>�?            �B@������������������������       ��r����?             >@������������������������       �؇���X�?             @������������������������       �                     @        #                   �^@�LQ�1	�?             G@!       "                    �?�eP*L��?             &@������������������������       �                     @������������������������       �      �?              @$       %                   `^@��?^�k�?            �A@������������������������       �                     �?������������������������       �                     A@'       ,                    �?�:�]��?�            �i@(       +                    �?�nkK�?r             g@)       *                    c@Х-��ٹ?]            �b@������������������������       �/\a��?V            �a@������������������������       ��q�q�?             "@������������������������       �                     A@-       0                   �q@���Q��?             4@.       /                    @z�G�z�?             .@������������������������       �և���X�?             @������������������������       �                      @������������������������       �                     @�t�bh�h(h+K ��h-��R�(KK1KK��ha�B        r@     pt@     �k@     �X@      E@      J@      3@      C@      *@              @      C@             �@@      @      @      7@      ,@      5@      @      0@      @      @               @      "@              @       @      @     �f@     �G@     �f@      E@     �L@      A@      <@      =@      =@      @     �^@       @     �^@      @               @              @     �P@     �l@      I@      D@      $@      A@      $@      ;@      @      :@      @      �?              @      D@      @      @      @      @              @      @      A@      �?              �?      A@              0@     �g@       @      f@       @     �a@      @      a@      @      @              A@       @      (@      @      (@      @      @               @      @        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ�]_AhG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK3hyh(h+K ��h-��R�(KK3��h��B(                             �?�:�Ӛ��?�           8�@              
             �?^���u��?�            pp@       
       	          pff�?�����?t             e@                           �?`՟�G��?             ?@              	          833�?"pc�
�?             &@������������������������       �                      @������������������������       �                     "@       	       	          833�?      �?             4@������������������������       �$�q-�?
             *@������������������������       �և���X�?             @                           @ ���v�?^             a@                            G@���7�?             F@������������������������       �z�G�z�?             @������������������������       � ���J��?            �C@������������������������       �        A            @W@                           �?�o+��?@            �W@                          �d@��S�ۿ?             >@������������������������       �                     :@                           �?      �?             @������������������������       �                      @������������������������       �                      @              	          ��� @�n_Y�K�?,            @P@              	          ����?��~R���?+            �O@������������������������       �<|ۤ$�?&            �K@������������������������       �                      @������������������������       �                      @       &                   �l@�7�A�?�             v@       !       	          ����?�����?X            �b@                           �?�����?Q             a@������������������������       �                     J@                            �?h�����?5             U@������������������������       ���2(&�?             6@������������������������       �        &             O@"       %                   ``@�8��8��?             (@#       $                    �F@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @'       ,                    �?*Mp����?t            �i@(       )                   �m@���;QU�?-            @R@������������������������       �                      @*       +                    �?0z�(>��?,            �Q@������������������������       �        "            �L@������������������������       �d}h���?
             ,@-       0                   e@���˅��?G            ``@.       /                    @�q�q�?0            �V@������������������������       �      �?             <@������������������������       �r֛w���?             O@1       2                    �?,���i�?            �D@������������������������       ��?�|�?            �B@������������������������       �                     @�t�bh�h(h+K ��h-��R�(KK3KK��ha�B0       `q@     u@     @h@     @Q@      c@      0@      1@      ,@       @      "@       @                      "@      .@      @      (@      �?      @      @     �`@       @      E@       @      @      �?      C@      �?     @W@              E@     �J@       @      <@              :@       @       @       @                       @      D@      9@      D@      7@      @@      7@       @                       @      U@     �p@      ,@     �`@      @     �`@              J@      @     @T@      @      3@              O@      &@      �?      @      �?              �?      @               @             �Q@     �`@      @      Q@       @              @      Q@             �L@      @      &@     @P@     �P@      N@      >@      ,@      ,@      G@      0@      @      B@      �?      B@      @        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJL�OhG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK9hyh(h+K ��h-��R�(KK9��h��Bx                             �?b�#�(��?�           8�@                           @L@��3Fi�?            y@       
                    @(޻��?�            `l@                           �?�~
	�?z            �f@                           �? ���J��?g            �c@������������������������       �        <            @V@������������������������       ��L#���?+            �P@       	                   �\@H%u��?             9@������������������������       �      �?             @������������������������       �                     3@                           �?nM`����?             G@                          xp@���@��?            �B@������������������������       �����X�?             <@������������������������       �                     "@������������������������       �                     "@                           @r�%���?v            �e@                           @O@.��Zr��?C            @X@                           �?~|z����?%            �J@������������������������       ����"͏�?            �B@������������������������       �        
             0@                           �?��2(&�?             F@������������������������       �                    �@@������������������������       ��eP*L��?
             &@                          �d@�99lMt�?3            �S@                           b@8����?,            @Q@������������������������       �                     @������������������������       ���&����?*            @P@                          pq@�<ݚ�?             "@������������������������       �                     @������������������������       �                      @       ,       
             �?�(� ��?�            �j@        '       	          ����?��[�m�?c            �c@!       $                    �?     8�?'             P@"       #                   @]@d��0u��?             >@������������������������       �                     "@������������������������       ��G��l��?             5@%       &                    �N@�IєX�?             A@������������������������       �                     ;@������������������������       �����X�?             @(       +                    �?`�q�0ܴ?<            �W@)       *                    @�NW���?#            �J@������������������������       �`2U0*��?              I@������������������������       ��q�q�?             @������������������������       �                    �D@-       4                    @P@ؓ��M{�?            �K@.       1                   0n@D�n�3�?             C@/       0                   @j@����X�?             5@������������������������       ����Q��?             $@������������������������       �                     &@2       3                    @j���� �?             1@������������������������       �                     @������������������������       �                     $@5       6                    ]@�t����?             1@������������������������       �                     &@7       8                   �q@�q�q�?             @������������������������       �                      @������������������������       �                     @�t�bh�h(h+K ��h-��R�(KK9KK��ha�B�       �q@     �t@     @]@     �q@      B@     �g@      @     �e@      @      c@             @V@      @     �O@      @      6@      @      @              3@      =@      1@      =@       @      4@       @      "@                      "@     @T@     �W@      ?@     �P@      9@      <@      "@      <@      0@              @      C@             �@@      @      @      I@      <@      H@      5@              @      H@      1@       @      @              @       @             �d@     �H@     �`@      9@     �E@      5@      &@      3@              "@      &@      $@      @@       @      ;@              @       @     �V@      @     �H@      @      H@       @      �?       @     �D@              ?@      8@      0@      6@      @      .@      @      @              &@      $@      @              @      $@              .@       @      &@              @       @               @      @        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ��lhG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK+hyh(h+K ��h-��R�(KK+��h��Bh	                            pb@�FF,���?�           8�@              	          pff�?��X��?�            �q@                          @[@      �?3             U@������������������������       �                     ,@              	          pff�?�z�G��?+            �Q@                           �J@֭��F?�?            �G@������������������������       ��X�<ݺ?
             2@������������������������       ��f7�z�?             =@	       
                    �?�LQ�1	�?             7@������������������������       �                     0@������������������������       �և���X�?             @                          @\@(1�Fh�?�            �h@                           @Q@8�A�0��?             6@                          �l@�����?             3@������������������������       �      �?              @������������������������       �                     &@������������������������       �                     @                           @ܷ��?��?r            �e@                           �?�����D�?(            @P@������������������������       �Du9iH��?            �E@������������������������       �8�A�0��?             6@                          �e@��Ujѡ�?J            @[@������������������������       �P�c0"�?G            @Z@������������������������       �                     @       (       	          ���@����s��?�            �t@       !                    @�z�G��?�             t@              	          033�?P���Q�?�             n@                           c@@�R��?�             m@������������������������       ��{3/o"�?�            �k@������������������������       ��z�G��?             $@                            �?����X�?             @������������������������       �                      @������������������������       �                     @"       %                   �n@R�����?0             T@#       $                    �?Dc}h��?"             L@������������������������       ��KM�]�?             C@������������������������       ��E��ӭ�?             2@&       '                    �?r�q��?             8@������������������������       �      �?              @������������������������       ���2(&�?             6@)       *                    �H@��S�ۿ?
             .@������������������������       �                     �?������������������������       �        	             ,@�t�bh�h(h+K ��h-��R�(KK+KK��ha�B�       �o@     �v@     �g@     �V@      5@     �O@              ,@      5@     �H@      2@      =@      �?      1@      1@      (@      @      4@              0@      @      @      e@      ;@      *@      "@      *@      @       @      @      &@                      @     �c@      2@     �J@      (@      D@      @      *@      "@     �Y@      @     �Y@       @              @     �O@      q@     �H@     �p@      (@     �l@      $@     �k@      @      k@      @      @       @      @       @                      @     �B@     �E@      1@     �C@      @      A@      *@      @      4@      @      �?      �?      3@      @      ,@      �?              �?      ,@        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ�-#hG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK1hyh(h+K ��h-��R�(KK1��h��B�
                             �?�>$�*��?|           8�@                           �?v ��?�            �r@       
                    �?��d��?[            �d@                           @T�iA�?(            �Q@                            N@ףp=
�?             >@������������������������       �                     6@������������������������       �      �?              @       	                    \@P���Q�?             D@������������������������       ����Q��?             @������������������������       �                    �A@                          �b@��E�B��?3            �W@������������������������       �                     C@                          pc@d}h���?$             L@������������������������       ��q�q�?             .@������������������������       �������?            �D@              	          033�?�v��\�?\             a@                           �?�n_Y�K�?,            @P@                          �b@���j��?             G@������������������������       ����N8�?             5@������������������������       ��q�����?             9@                           �?p�ݯ��?             3@������������������������       �      �?              @������������������������       ��C��2(�?             &@              
             �?�X�<ݺ?0             R@������������������������       �        )             N@                           @�q�q�?             (@������������������������       ������H�?             "@������������������������       �                     @       *       	          033�?�Z;EF�?�            �s@       #                   �^@jO�9���?�            @o@       "                    @�:nR&y�??            �W@        !       	          ����? rpa�?>            @W@������������������������       � ��PUp�?.            �Q@������������������������       �"pc�
�?             6@������������������������       �                      @$       '                    �?�4�����?^            `c@%       &                    �?�S����?>            �W@������������������������       �                     A@������������������������       ��jTM��?&            �N@(       )       	          ����?�q�q�?              N@������������������������       �~�4_�g�?             F@������������������������       �                     0@+       0       
             �?     ��?(             P@,       /                    �?�^����?&            �M@-       .                   0b@�q�q�?             5@������������������������       ��<ݚ�?             2@������������������������       �                     @������������������������       �                     C@������������������������       �                     @�t�bh�h(h+K ��h-��R�(KK1KK��ha�B       �p@     �u@      d@     �a@     �J@     �[@     �D@      =@      @      ;@              6@      @      @      C@       @      @       @     �A@              (@     �T@              C@      (@      F@      $@      @       @     �C@      [@      =@      D@      9@     �@@      *@      4@      �?      *@      (@      @      (@      @       @      �?      $@      Q@      @      N@               @      @       @      �?              @     @[@     �i@     �L@      h@      @      V@      @      V@      �?     �Q@      @      2@       @              I@     @Z@      .@      T@              A@      .@      G@     �A@      9@      3@      9@      0@              J@      (@      J@      @      ,@      @      ,@      @              @      C@                      @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ5�;5hG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK+hyh(h+K ��h-��R�(KK+��h��Bh	                             �?����/��?�           8�@                           �?�b��-8�?�            �s@              
             �?\������?N            �[@������������������������       �                     5@                           @����E��?@            �V@                          �]@�z�G��?*             N@������������������������       �                     @������������������������       ��<ݚ�?'             K@	       
                    �?�������?             >@������������������������       ��KM�]�?             3@������������������������       ��eP*L��?	             &@              	          033�?�d2 Λ�?�            �i@                           @M@���L��?u            �f@                           �?`�q�0ܴ?[            �a@������������������������       �        (            �M@������������������������       ���p\�?3            �T@                          �p@�p ��?            �D@������������������������       �                     <@������������������������       ���
ц��?             *@                           �?      �?             6@                          �h@�n_Y�K�?	             *@������������������������       �                     @������������������������       �z�G�z�?             $@                          �^@�q�q�?             "@������������������������       �                      @������������������������       �؇���X�?             @                           �E@V��~��?�            �r@������������������������       �        	             *@       $                    @��r._�?�            �q@       !       
             �?�,A7H�?U            ``@               
             �?��Lɿ��?3            �T@������������������������       �     ��?	             0@������������������������       ��L#���?*            �P@"       #                    �?r�q��?"             H@������������������������       ��z�G��?             >@������������������������       ��E��ӭ�?             2@%       (                   �a@ȵHPS!�?[            �c@&       '                    �?���(-�?/            @R@������������������������       �                     ?@������������������������       �@4և���?             E@)       *                    �?b:�&���?,            �T@������������������������       �@��8��?             H@������������������������       ����Q��?            �A@�t�bh�h(h+K ��h-��R�(KK+KK��ha�B�       0t@     @r@     @U@     �l@      O@     �H@      5@             �D@     �H@      2@      E@      @              (@      E@      7@      @      1@       @      @      @      7@     �f@      (@     @e@      @     �`@             �M@      @      S@      @     �A@              <@      @      @      &@      &@      @       @      @               @       @      @      @               @      @      �?     �m@      O@              *@     �m@     �H@      Y@      ?@     �R@      "@      &@      @     �O@      @      :@      6@      5@      "@      @      *@     @a@      2@     �Q@      @      ?@             �C@      @      Q@      .@     �G@      �?      5@      ,@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJi4�hG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK5hyh(h+K ��h-��R�(KK5��h��B�                             �?8�! ���?�           8�@                           �?��ܭ��?�            s@       
                    @��E�@�?\             b@                           �?���O1��?5            �T@                          �\@���Q��?             @������������������������       �                      @������������������������       ��q�q�?             @       	                    �?�ݜ�?1            �S@������������������������       ���ϭ�*�?&             M@������������������������       �      �?             4@              
             �?`��:�?'            �N@                          �c@ qP��B�?            �E@������������������������       �                     C@������������������������       �z�G�z�?             @                           �?b�2�tk�?
             2@������������������������       �r�q��?             @������������������������       �r�q��?             (@                          Xp@��	l�?i             d@                           @���E�?9            �U@������������������������       �                     8@                          @[@ ������?*            �O@������������������������       ��q�q�?             @������������������������       �        '             N@                           �?������?0            �R@                          @`@X�<ݚ�?             2@������������������������       ����!pc�?             &@������������������������       �                     @������������������������       �        $             L@       ,       
             �?��a�n`�?�            `s@       %       	          033�?\X��t�?N            �\@       "                    @l��
I��?5            @T@        !                    �?�����?             E@������������������������       �                     =@������������������������       ��	j*D�?             *@#       $                   �_@Hث3���?            �C@������������������������       �8����?             7@������������������������       �     ��?
             0@&       )                    `@������?             A@'       (                   �j@�IєX�?             1@������������������������       �      �?             @������������������������       �                     *@*       +                    �N@j���� �?             1@������������������������       ��<ݚ�?             "@������������������������       �      �?              @-       4       	          hff@��-�=��?w            `h@.       1                   c@��8���?u             h@/       0                    �?��V#�?             �E@������������������������       ��LQ�1	�?             7@������������������������       ��G�z��?             4@2       3                   �c@�'F�3�?U            �b@������������������������       ��LQ�1	�?             7@������������������������       �        H            �_@������������������������       �                     @�t�bh�h(h+K ��h-��R�(KK5KK��ha�BP       �q@     �t@     �j@      W@     �N@     �T@      (@     �Q@       @      @               @       @      �?      $@      Q@      @     �J@      @      .@     �H@      (@      E@      �?      C@              @      �?      @      &@      @      �?       @      $@      c@      "@     �U@      �?      8@              O@      �?       @      �?      N@             �P@       @      $@       @      @       @      @              L@             �Q@      n@      I@     @P@      8@     �L@      @      C@              =@      @      "@      4@      3@      @      0@      *@      @      :@       @      0@      �?      @      �?      *@              $@      @      @       @      @      @      4@     �e@      1@     �e@      ,@      =@      @      4@      &@      "@      @     @b@      @      4@             �_@      @        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ�ThG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK+hyh(h+K ��h-��R�(KK+��h��Bh	                             @D^��#��?�           8�@              	          `ff @� u��?�            �u@       
                    �?r�'�Z�?�            �s@                           @M@���;QU�?�            `k@                          `_@�Sa��?n            �d@������������������������       �"pc�
�?	             &@������������������������       �@f����?e            �c@       	       	          ����?�θ�?"             J@������������������������       �$��m��?             :@������������������������       �ȵHPS!�?             :@                           �?ڡR����?>            �X@                           �? ���J��?            �C@������������������������       �                     ?@������������������������       �      �?              @                           �?L
�q��?%            �M@������������������������       ���r._�?            �D@������������������������       ��E��ӭ�?
             2@                           \@д>��C�?             =@������������������������       �                      @                           �?�����H�?             ;@              
             �?�z�G��?             $@������������������������       �      �?             @������������������������       �                     @������������������������       �                     1@                          @[@0�".���?�            �p@                           Y@������?
             1@                          `c@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     (@       $                    �?�9���[�?�            �o@        !                    �?��(!i�?x            �h@������������������������       �        >             W@"       #                    �L@B�����?:             Z@������������������������       ���v$���?#            �N@������������������������       ��K��&�?            �E@%       (                   �l@h�����?#             L@&       '       	          `ff�?���Q��?             9@������������������������       ��q�q�?	             .@������������������������       �                     $@)       *                   �\@�4�����?             ?@������������������������       �                      @������������������������       ��c�Α�?             =@�t�bh�h(h+K ��h-��R�(KK+KK��ha�B�       �q@     �t@     �S@     �p@     �K@     `p@      .@     �i@      @     �d@       @      "@      �?     `c@      (@      D@      "@      1@      @      7@      D@      M@      �?      C@              ?@      �?      @     �C@      4@      A@      @      @      *@      8@      @               @      8@      @      @      @      �?      @      @              1@             �i@     �O@      @      *@      @      �?              �?      @                      (@     @i@      I@      f@      3@      W@             @U@      3@      N@      �?      9@      2@      9@      ?@      .@      $@      @      $@      $@              $@      5@       @               @      5@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ5�R/hG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK7hyh(h+K ��h-��R�(KK7��h��B                             @K@r � 	��?�           8�@                           @0էu���?�            �r@              	          033�?������?            �i@                           ^@���g�?u            �g@������������������������       �                     @              	          ����?@�Gpm��?q             g@������������������������       �h㱪��?A            �[@������������������������       �        0            �R@	       
                    �?����X�?
             ,@������������������������       �                     @              	          ���@X�<ݚ�?             "@������������������������       �                     @������������������������       �                     @                           �?(���@��?@            �W@                          �a@D7�J��?#            �K@������������������������       �                     &@                          Pd@���|���?             F@������������������������       �        
             2@������������������������       ��n_Y�K�?             :@                          �e@�7��?            �C@              
             �?�?�|�?            �B@������������������������       �                     =@������������������������       �      �?              @              	          ���@      �?              @������������������������       �                     �?������������������������       �                     �?       *       	          033�?�,�٧��?�            �s@       #                    �?�JS���?�            �k@                            �?�e0����?X            �a@                           @��k��?$            �J@������������������������       ����B���?             :@������������������������       ������H�?             ;@!       "                    �?�<ݚ�?4            �V@������������������������       ���V#�?            �E@������������������������       ���E�B��?            �G@$       '                    �?��Sݭg�?-            �S@%       &                    �?�nkK�?             G@������������������������       �����X�?             @������������������������       �                    �C@(       )       	          ����?     ��?             @@������������������������       �z�G�z�?             4@������������������������       �r�q��?             (@+       0                   �a@�KM�]�?>            �W@,       /                    @���U�?%            �L@-       .                    �?���}<S�?             7@������������������������       �                     *@������������������������       �z�G�z�?             $@������������������������       �                     A@1       4                    @���y4F�?             C@2       3                    �?`Jj��?             ?@������������������������       �                     <@������������������������       ��q�q�?             @5       6                   b@؇���X�?             @������������������������       �                     �?������������������������       �r�q��?             @�t�bh�h(h+K ��h-��R�(KK7KK��ha�Bp       @q@     0u@      U@     �j@      4@      g@      $@     �f@      @              @     �f@      @     �Z@             �R@      $@      @      @              @      @              @      @              P@      >@      ;@      <@      &@              0@      <@              2@      0@      $@     �B@       @      B@      �?      =@              @      �?      �?      �?              �?      �?              h@      _@     �Z@     �\@     �H@     �W@      =@      8@      @      5@      8@      @      4@     �Q@      ,@      =@      @     �D@      M@      4@      F@       @      @       @     �C@              ,@      2@      @      0@      $@       @     @U@      $@     �K@       @      5@       @      *@               @       @      A@              >@       @      =@       @      <@              �?       @      �?      @              �?      �?      @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ�%hG        hNhG        hGKhHKhIh(h+K ��h-��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh(h+K ��h-��R�(KK��hP�C       �t�bK��R�}�(hKhxK7hyh(h+K ��h-��R�(KK7��h��B                             �?���i��?�           8�@                           �?��hY��?�            r@       
                     N@     ��?R             `@                           @L@��j2��?@            @Y@              
             �?��=A��?4             S@������������������������       � s�n_Y�?#             J@������������������������       �r�q��?             8@       	                   `a@z�G�z�?             9@������������������������       �                     4@������������������������       �                     @                          P`@�+$�jP�?             ;@                           �Q@�q�q�?             "@������������������������       �                     @������������������������       �                     @                          `g@�����H�?             2@������������������������       �                     �?������������������������       ��IєX�?             1@              	          ����?���`uӽ?l             d@                           @������?             A@                          �_@      �?             0@������������������������       �r�q��?
             (@������������������������       �                     @                           @O@�����H�?             2@������������������������       ��IєX�?             1@������������������������       �                     �?                           �O@ ���z��?S            �_@������������������������       �        B             X@                            P@`Jj��?             ?@������������������������       ��q�q�?             @������������������������       �                     <@       .                   �a@v�PT!�?�            `t@        '                   Pa@��S���?(             N@!       $       	          `ff�?���"͏�?            �B@"       #                    `@ףp=
�?             >@������������������������       �d}h���?             ,@������������������������       �        	             0@%       &                    @P@؇���X�?             @������������������������       �                     @������������������������       �                     �?(       +                   �a@�㙢�c�?             7@)       *                    �?      �?	             0@������������������������       �                     �?������������������������       ���S�ۿ?             .@,       -                    �?����X�?             @������������������������       �                      @������������������������       �                     @/       0                    �?���܉Z�?�            �p@������������������������       �        @            @Z@1       4                    @L@���z��?j             d@2       3       	          `ff@����&��?D            �Z@������������������������       ��b�E�V�?A            �Y@������������������������       �                     @5       6                    �?\�����?&            �K@������������������������       �k��9�?             �F@������������������������       ��z�G��?             $@�t�bh�h(h+K ��h-��R�(KK7KK��ha�Bp       0r@     @t@     �k@     �P@      R@      L@      I@     �I@     �F@      ?@     �D@      &@      @      4@      @      4@              4@      @              6@      @      @      @      @                      @      0@       @              �?      0@      �?     �b@      $@      :@       @      $@      @      $@       @              @      0@       @      0@      �?              �?     @_@       @      X@              =@       @      �?       @      <@              Q@      p@      <@      @@      "@      <@      @      ;@      @      &@              0@      @      �?      @                      �?      3@      @      ,@       @              �?      ,@      �?      @       @               @      @              D@     @l@             @Z@      D@     @^@      &@     �W@       @     �W@      @              =@      :@      :@      3@      @      @�t�bubhhube�oob_decision_function_�h(h+K ��h-��R�(KMgK��ha�Bp&  w��zNu�?p̥0V1�?N�{��?A��Ѐ��?�x#�?z��>��?n���?�H��=�?�0�&�?�=��d�?C>gm���?p0�$HL�?%܃T��?j�𕯚�?
k1���?�)��"��?m�wܷ?@q}�?����q��?E�zp�?�.s͸?#��Q��?���>�?�/�@L�?�NKx��?#K�~h�?�E���?��{_���?�MR����?O���O(�?�cV��_�?�3�-��?�m��A�?�#\�ŗ?�)�0ƫ?h�%��C�?!Py`��?�_?K��?<h9�
�?���q\=�?�;3���?%!f��R�?�ŷA���?Cɗ��?0yWJ?��?8D�(�?�┽ͷ?��cMH�?1�qZ�?�;�;��?C��+�?^,sjp�?Ð�)�ը?�&`��r�?��I9D�?�8[c���?h~:4��?�\,^F�?�	}�e�?H���Ѵ?q'$0���?G��率�?]�ڢ3�?�v��.f�?
��)�~�?|�@�?�S��E��?�u�F׏�?!�����?�r&)��?�I�&��?����ek�?	��[�1�?�#�r�?�GDʋ�?���[C��?{W����?AT}���? $�%���?��
��?�42#�?0���Ν�?�w���?7���W~�?�Y#�$��?˔�o۫�?~���vֻ?��&1��?N���߯�?�5���?�������?�ݏ����?�E�7���?�t���Z�?K��|���?,�1���?^�ߥB�?G�@�z��?E��I/ם?eZ��F�?^+��3�?��n�c�?O`����?�O����?q�)���?F��9��?vI����?�mgjL�?bӅn 	�?O��o��?B��B��?^��^x
�?sο���?���,�?�������?��J���?���kv�?�}����?� d�{��?��oZj�?H �YYz�?�S�B�?�ih�?�?�l��?��W�s1�?�2Fg�?�Y	�s��?�����?P+����?b��H<��?�{�Ev�?���B7��?�4��ߙ�?�,|���?����=�?%�	r2a�?H3_�ȱ?��t���?\𷴍p�?�Ғ���?�HL�\��?���(��?+Aa�0��?�}=o�}�?�����?��ub�?-;�&N��?�&�ʎ=�?��E���?H]IWh��?fh��ߥ�?ȼc Ѻ?�;Ɖ��? #6ϱӲ?^���BM�?���+�?��>?���?�+����?��;}��?� f�?����-��?�*��޳?"�(l+�?��Ij��?6^��I#�?�P>,[��?1���?�����?�}�z�?�]��Ua�?�	�~�?�^�>p�?Ҙ�I�?c9뱽��?��!�9a�?�3�0��?ΣĪ�?b�v����?�g�,�?��ɐ>��?�a�p%��?!��{�>�?�qN7��?vq�E�ٷ?���2�:�?.��ٮ8�?�w����?�|D���?*�.mS�?l�-ɪ�?�}��?OF����?���Y.��?B��0���?��X�]��?���њ�?%O�/oA�?gҗ?��G|0�?0~(����?�2� M9�?���[֘�?y�Յ2��?=LR�k&�?�����C�?�x�� ��?b��B�/�?�/����?�u�s��?5�k�?�yG���?��!�|�?9�U6�?����U��?����2<�?�8�5�?�{4aP��?�"\�|��?@�)g��?p��5�?�����?��-�w�?�J [�!�?���o�?ר��e��?��C�`�?\��`W��?���'��?�T	��/�?Ԫ}���?�CQ<�&�?^����?:p���e�?�#����?d|���R�?<�$q�z�?ɹ��?n�0����?X0�9��?�>�K_�?[�l�6��?ӕɪ��?Ϭҷ��?��T��?��5��m�? e���?�>�Z;�?ςqJ���?3\�-.�?�Q����?���?@x�?G�q�=�?/��˯�?��Ih��?�un ��?�(F~�K�?G�,��?���?��?���rE�?�s
u�?����Z��?����R��?F��4�)�?�]yYβ�?�bJ�
�?�tֲ ��?���Jb$�?㢶s;�?�������?�>�����?tD�_!��?���wS�?� dc��?���3n�?f��)v��?�P�u���?�+;�i�?�)j�$K�?:��Je�?l�1V���?HƼ\��?�6ghTE�?~��Tw�?���UD�?�A��QU�?=��pU�?�w.ݮΡ?�-��?^�l�?@�?or��?�D�����?�]��*�?rx����?aD���?�"���? ~�� ��?o��#1��?�+n�-�?��@�[�?�3����?�DR���?��V�/��?l�
֗?�4?�OA�?,�8�#��?�嘌�O�?��"Q�m�?��nW��?���t��?2
=lѫ�?��G0�?+ �����?C=�I���?}��l�~�?���{���?���]�?�NM ��?��%���?�+O9��?�Gk�ӯ?k��o��?I��y�?8��
�?>D�R�~�?�`4��?󹌿~F�?^]g��,�?*�ɧ5��?b�9����?��I�?��?1���?�:���"�?$�޸w�?ʷ�B��?��l�7�?�C��2�?D�ƫE�?w?�s�t�?!�'/#�?{�cCs�?�]mu��?�'*����?��te�3�?�efQӌ�?���P��??�
�k��?��@���?�/���?��D��?ײ�r�?�D���?�݈��$�?�t�#���?�"�Ղ�?�BDOe�?ջ����?h��0��?L�����?x誦���?G��ʒ��?��c�C�?��G�3��?�j��E��?�J�6݉�?������?���;���?u��h�?rš��K�?���.��?Xh;�Fj�?V��mV�?wȐdO5�?��v�?�?<@B-��?!(��)��?�}��e=�?H�z�y�?m'�
=�?��/
�e�?�)�z&��?��恊��?WZ�_�L�?�G�6��?�^�둜�?���~��?M���?�ΓT��?�ö
��?����?'$>�#�?u7Û��?
��C��?���<���?@$�a6��?JC����?,�ߕ���?_0���?�g����?
��cG��?`É���?��C�.�?0���(��? ����?�o��!�?/�佊�?h7����?u�Ş���?]l�	S�?�K���???����?�F�����?p�~�U��?�����?��}!D�?G�>d��?sc�7��?.�����?A/���;�?n^Ӗ5v�?3�%M9��?xh\�E�?���Q��?+�
����?Oկ%��?˯��Z��?�� �?�ϛ}��?CV.�?X��a��?����)/�?�xg޿9�?�C� ��?�c�����?e���Q��?Iк��?�})�8"�?ń�-*y�?�=�j��?��_�NH�?�0����?��+%�?B�N����?��zԥ�?�	����?�l��O�?j�\A_��?�P+ŭ��?��ZG�h�?@+.�ta�?����X��?��A�/9�?��|����?�9�7׳?c�X��?uV�6d�?�T�����?���z�;�?3*n
y��?1�����?vWP�8�?�e�4#��?�f�2���?T�#����?�:�����?��+�c��?������?c���?8�3����?�n��?�t�ȍ��?�s��?�?c�pz�?�j��8�?��<���?��3��?�d?�?C��w�?J�RD�?Sh(�Ϧ�?h��&�ɲ?^b�Œ�?P���6�?S��a���?r���?�/�?��;=4�?�Y���?�d�uϯ�?/¿^���?��
ʲ?���Ӳ �?1A���?�i�}���?�A%1�?�|�C4/�?�`�24�?�7?ssi�?�-�?C}�����?��2�?����o�?<��?
��x���?{���3 �?���"�g�?����[�?uHL�;T�?(��v��?]AP�?�E�}_��?J�>?=Ǵ?8$Xg�?C��Z{�?�+1RJخ?��C����?��QQ��?�Sޡ��?���7�?@N�E`��?p���g�?���6{8�?�d$��8�?3�
o!�?7/�C�{�?���N��?���r��?C���F�?�^R��?�%�#��?�n�v�?��e���?W�����?��x(��?���5��?�﵊|�?��@(��?��AV�?0�r����?:'G��?����6?�?g�%!�P�?�)��M��?e�M��?j�Ȫ���?�%��>�?�v��Op�?C�g�̴�?|{0�f��?����y�?pM Ͱ��?��ĭv}�?_ǎT���?K�ێݒ�?[�8�6�?���z���?�� ��?<�n9�?'�4&�?�i�D��?K�]9�?��6�fC�?.�d�L^�?{�2!Xa�?����ԓ?�Pg��?��usK�?�b�K�?��N�Z�?�a��N,�?�s!v��?�Y��fy�?�3�(�4�?��J�ai�?f!���Ӓ?����X0�?����9�?�)P��?���v2�?���BX�?�[V>zO�?��k�?�?>�T��?�-��8��?�t�q��?x9����?Ә��`�?;�jj���?�*+u.�?��}����?��0���?=�f�m�?�.,��'�?C;7i�9�?��r���?eTh���?��eW��?:�=$L�?�Bx;|��?�Aߢ�?����?��`F���?���{Pd�?�sߏ��?��7�?��N ޸�?"���#�?Ĭ7kH��?w��)o�?�h�D�!�?�e�n�7�?e�/��?��$��c�?������?���mV�?\�m����?F�$�2�?	y��?����7�?H>MHP'�?m���+��?��Fx���?��=d*�?��k��?y.J'|�?m��D&k�?�*h7�r�?S$��?��ێ��?�1����?f����T�?�gyN��?L�����?��*ۊ�?��S�&��?�+�_e�?��Sǁj�?䤨���?��+��s�?�V��$\�?lK=���?��N�u��?�%N���?�ʥԗ)�?R���f�?������?����M��?ޱf�/S�?E�2�Y�?=��9�?�'��Q��?}�L!*�?!�w5�?��
il��?.��rr+�?Cm�	�?�%�	���?�έRH�?M�T+�-�?�Rb)�?Zk罵;�?��hô��?��K�%��?H�tNz��?ղ-���?5~���y�?X9��jĐ?���m�m�?*�F2Or�?ǿ�~��?� a,�?�������?�?3��?:T�NG��?�սXܫ�?����{�?B��@8�?�7c�o��?B�|���?=�+npٽ?��:��D�?	�$)5Ȧ?p�m�|��?<٦|.�?�I��`t�?sߏ�4��?d��Yf�?B5���?���*#�?�����?���- �?�ա��?��{��? �'ݺ�?�k`ˋ�?8	��p�?=o�����?��S]A	�?&�U����?V�wV�?��8bj��?
���c��?z�*0N �?��8R��?���֍��?R*+,�?W�j����?S��N��?�"v�}�?��ˎo��?�s���|�?u�p|;�?Y,z$�?��Ə���?6�Ɂ{�?�yڥ��?fbh^�U�?�<'���?�vO�C�?�1�Ă�?����v��?�j�����?�ʵ�?�dy�O�?ʦ!�>��?��tU��?���/���?���~�_�?8$�x�?����N�?, c�/$�?@�Ⱥ�? �_���?$�_�&��?� 
���?];��4��?'��YNB�?V�XI�t�?ԮS[�E�?��afv�?(*<3��?lK,?z�?&�4p���?�#�k��?������?�o&s��?z��fD��?\�́��?�b ����?�?o�f�?�;0$Q��?���-��?���H��?�m|�y��?��"Î�?��0��?�~��~�?lw���?N"�! �?J���q�?j��,��?�`�9l��?���Ʌ�?F��L��?ܼr�ك�?5�����?�s?(��?��,��(�?��t����?�~J�u��?��(��?�xK��[�?fi}�H�?i�E�?�-�t���?#��7�\�?t�!���?�}�$��? h�ݐQ�?�n���O�?e"��`�?^g%�:�?)�6Kqy�?{��oT��?"�
�*��?��5�n�?bF�� 2�?5��)�?�k�^���?��r_�I�?��4�f��?��Uf��?h@5SJ��?-C�+��?�4��:��?��D����?���lT�?��	s�?�oϸ��?��c�+�?�N<����?@X/7���?�O�����?ZP����?�� �q<�?Bt�S0��?���?+���a��?N��ux��?���+�?.��8���?��2w�?yEH�;b�?��i���?�B�l� �?�Y?�?�?�1�� �?h`�% �?�ϐy�o�?Y��յ?ߔC�AE�?W}�Q��?,��J���?�L���?4�g�� �?R�3Aȳ?7������?Y��1�?T�!�|g�??��"���?�AK�U��?;N�0t�?#���^�?�Zg�Q�?*�b�? �J���?��Z���?0)�E |�?�ZB�{��?�5f�Ϻ?C9s���?����`�?�É����?]9�hbP�?�����?SR$j�?�Y�[�+�?[���5��?�-BAY)�?�z�O�?�����?.O\�U��?v�DU �?xڰ���?W�4?g�?������?�я�L�?̨�` �?�2����?L�];w�?UM��#�?Pm�l6`�?�JzL&�?�d?7�?l��#�?Y���\��?��A�F�?I�f�w�?~o���?��.%�#�?�������?T='��?�W�ٱ��?�[�7#��?�2���?���I��?�#���?)��U��?�cNT���?l�K����?��v�`��?�_
1 t�?��w�^�?��쯿�?�c�M@�?l_����?JP<*��?�|�%��? ࠕ���?�S�?�?����8�?U�t����?W�E��?�;��&�?�8O'[b�?�m1u���?GH:+j	�?����V�?֢��$#�?=m`���?.����>�?uZ��?�҄�<��?O�B<n�?�
��G�?=��&g�?Y�!�?gf k�a�?33�)A<�?߬�Z�P�?���ҫ��?(W���?�k�r�?//�s���?�����?9xAY�?��}M�?�f����?�L�~;��?���в}�?ㄶ��$�? �@N0�?B�o~�3�?VS��?{�oOeU�?7�hO���?M���}�?��+0�?��u�g�?�H`6��?p�~&���?�8�Ƙ�?\O���?�K���
�?-PH��?S�����?�:Y
�?v��}�6�?bʌ`X��?��a%,�?��O���?+�ri1�?<�G��3�?�\�A�?�wF-�|�?�Wg.6��?3:9��?��x��0�?$�Ö���?c?�0z<�?r�<�?q���{e�?ǀ�,B��?��9tk�?���x���?�������?��%���?�`IL��?c��͟-�?�؁�A�?*�N�l|�?i�Ԅc��?�����?E���$�?�"�m�?�*x�L�?��P"mv�?)��;D�?[L�pW�?5��H�?0x���?�����?h�l�_��?ť����?���yV��?���O�Z�?�kU�?�-�a3��?�1Of��?��˼�X�?��R;%�?W����??j�;��?���!&�?���坭?n�۴c��?��"Y�4�?����Y�?�����?k�a����?&�'Wђ�?�IY�˝�?�akZE#�?t-��i�?F�;0K��?�g\��?�vx�Q��?M�N�?�^.���?�H*ǮN�?�m5NTl�?C��F�&�?��"�,[�?�����?�| ��?��@�rP�?�D~{_�?S�ㄲ��?W/�����?�R��?����ݿ�?�}<Ц�?'/8���?]���U��?����?d� &4�?9}�����?� �P�?����^�?	�s�7��?~#r��?�y\�q��?�Go	�?Q���q�?sW.*��?C�pV��?��15g��?o_�t�?���h�?�������?P�ђ���?v�$'tu�?��6����?W�c�
��?�gD�	�?�Tz�D��?��B��"�?�� �t��?l���Y��?��d��?�<��7�?�0���?/���ˡ�?=fkϴ��?�LJ�%�?� 5+z�?g}+�S�?��;��?�\4/�?v��FX�?̆<���?�Л�^��?���м�?~|����?� �O�?�1���?p���GE�?0d��?��7E��?L�O����?k
lO��?H����7�?ܜ	���?;i�Qr�?my��x��?�0m�~�?��?KV�?� �l���?�?�d��?\'f�T��?�bg6���?�B0�+�?���s(j�?��K�?}G��}�?߮� ���?A�����?��7)ٮ?���lm�?�2/{@��?i�&��;�?�����?Q� �$�?��=.��?��G�;�?J,
��?j������?j�R+�?�W��S�?V�V��t�?Ա�,�E�?WU,I�?C�W�N��?��z� �?�^�0���?�7M��#�?G�,����? 6�#h�?���_�/�?�����?�rp>;�?',Qr�?fO���7�?��0{�K�?�<���?��
���?�DW���?����}�?�+#?N0�?��|z��?X7X�0�?�0�Xy�?��?��?�#t�H�?����o�?_9�6��?p5�K��?�*��r�?���F�?�{Y�ΰ?��4-��?�E��|��?��ݺt�?qPH�7K�?A��� ��?ܝ���T�?G�`x6V�?�G�ٿ�?�_�;f�?P��`<T�?敎�sx�?��y�9�?�[�3$1�?���$R�?��m���?��Z]��?�@{��S�?L�\|'�?Z��Ay��? �Lr~J�?�w�6��?3�k��?xfxʮ�?-���C7�?�-O���?j��(��?mI�vMΣ?x`�c: �?�s���;�?r<�>UA�?�q� X՗?a7�c�?�Df��?�o{��?B 	����?�޿j�{�?WP�	��?^�_CZ��?QP�Җ�?>��a�?��Da�?�4��?`��m���?#\,E�?w��i]��? �Յ�t�?��T���?�:�)Z¨?V<e]�s�?�[e��^�?�f�A(�?�_����? *�%o��?�Ѫ���?��]��2�?
�՚$�?bϣRv��?�J�h{�?_�rIX�?)�'�?���,���?��\�T�?n��>Z��?2��x�L�?�r�4[�?W�����?U���(��?o��i�?AB(��Y�?b�ҏe�?������?�B&�=�?t�;��?��Y��?��L���?��h݅�?��.�E��?k�����?�2H �?��u���?:�$	��?�m_{]��?��%e�?�춢��?���.�t�?LS��	��?<˪�a_�?#ō�O�?�\G�v�?'�6�ZV�?�����?�Z�C�1�?Pi���?�n"�.�?ٍ�O�?[��G�y�?�p��0�?ȧ��m�?�`�H��?� 6&�?����l��?�wsd-��?� 2nJ��?� ҭ��?�7o�±?���eIu�?���ѴU�?o�ʖ7~�?	)V���?�x^�µ�?��А��?�t�b�
oob_score_�hfhaC�\7�u��?���R�hhub.